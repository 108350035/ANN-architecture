module CHIP( 	
	// Inpt signals
	clk,
	rst_n,
	in_valid_d,
	in_valid_t,
	in_valid_w1,
	in_valid_w2,
	data_point,
	target,
	weight1,
	weight2,
	// Output signals
	out_valid,
	out
);
input  clk, rst_n, in_valid_d, in_valid_t, in_valid_w1, in_valid_w2;
input [31:0] data_point, target;
input [31:0] weight1, weight2;
output out_valid;
output  [31:0] out;

wire   C_clk;
wire   C_rst_n;
wire   C_in_valid_d,C_in_valid_t,C_in_valid_w1,C_in_valid_w2;
wire  [31:0] C_data_point,C_target,C_weight1,C_weight2;

wire  C_out_valid;
wire  [31:0] C_out;

wire BUF_clk;
CLKBUFX20 buf0(.A(C_clk),.Y(BUF_clk));

NN I_NN(
	.clk(BUF_clk),
	.rst_n(C_rst_n),
	.in_valid_d(C_in_valid_d),
	.in_valid_t(C_in_valid_t),
	.in_valid_w1(C_in_valid_w1),
	.in_valid_w2(C_in_valid_w2),
	.data_point(C_data_point),
	.target(C_target),
	.weight1(C_weight1),
	.weight2(C_weight2),
	.out_valid(C_out_valid),
	.out(C_out)
);

// Input Pads
PDUSDGZ I_CLK(.PAD(clk), .C(C_clk));
PDUSDGZ I_RESET(.PAD(rst_n), .C(C_rst_n));
PDUSDGZ I_IN_VALID_D(.PAD(in_valid_d), .C(C_in_valid_d));
PDUSDGZ I_IN_VALID_T(.PAD(in_valid_t), .C(C_in_valid_t));
PDUSDGZ I_IN_VALID_W1(.PAD(in_valid_w1), .C(C_in_valid_w1));
PDUSDGZ I_IN_VALID_W2(.PAD(in_valid_w2), .C(C_in_valid_w2));
PDUSDGZ I_D_P0  (.PAD(data_point[0]),  .C(C_data_point[0]));
PDUSDGZ I_D_P1  (.PAD(data_point[1]),  .C(C_data_point[1]));
PDUSDGZ I_D_P2  (.PAD(data_point[2]),  .C(C_data_point[2]));
PDUSDGZ I_D_P3  (.PAD(data_point[3]),  .C(C_data_point[3]));
PDUSDGZ I_D_P4  (.PAD(data_point[4]),  .C(C_data_point[4]));
PDUSDGZ I_D_P5  (.PAD(data_point[5]),  .C(C_data_point[5]));
PDUSDGZ I_D_P6  (.PAD(data_point[6]),  .C(C_data_point[6]));
PDUSDGZ I_D_P7  (.PAD(data_point[7]),  .C(C_data_point[7]));
PDUSDGZ I_D_P8  (.PAD(data_point[8]),  .C(C_data_point[8]));
PDUSDGZ I_D_P9  (.PAD(data_point[9]),  .C(C_data_point[9]));
PDUSDGZ I_D_P10 (.PAD(data_point[10]), .C(C_data_point[10]));
PDUSDGZ I_D_P11 (.PAD(data_point[11]), .C(C_data_point[11]));
PDUSDGZ I_D_P12 (.PAD(data_point[12]), .C(C_data_point[12]));
PDUSDGZ I_D_P13 (.PAD(data_point[13]), .C(C_data_point[13]));
PDUSDGZ I_D_P14 (.PAD(data_point[14]), .C(C_data_point[14]));
PDUSDGZ I_D_P15 (.PAD(data_point[15]), .C(C_data_point[15]));
PDUSDGZ I_D_P16 (.PAD(data_point[16]), .C(C_data_point[16]));
PDUSDGZ I_D_P17 (.PAD(data_point[17]), .C(C_data_point[17]));
PDUSDGZ I_D_P18 (.PAD(data_point[18]), .C(C_data_point[18]));
PDUSDGZ I_D_P19 (.PAD(data_point[19]), .C(C_data_point[19]));
PDUSDGZ I_D_P20 (.PAD(data_point[20]), .C(C_data_point[20]));
PDUSDGZ I_D_P21 (.PAD(data_point[21]), .C(C_data_point[21]));
PDUSDGZ I_D_P22 (.PAD(data_point[22]), .C(C_data_point[22]));
PDUSDGZ I_D_P23 (.PAD(data_point[23]), .C(C_data_point[23]));
PDUSDGZ I_D_P24 (.PAD(data_point[24]), .C(C_data_point[24]));
PDUSDGZ I_D_P25 (.PAD(data_point[25]), .C(C_data_point[25]));
PDUSDGZ I_D_P26 (.PAD(data_point[26]), .C(C_data_point[26]));
PDUSDGZ I_D_P27 (.PAD(data_point[27]), .C(C_data_point[27]));
PDUSDGZ I_D_P28 (.PAD(data_point[28]), .C(C_data_point[28]));
PDUSDGZ I_D_P29 (.PAD(data_point[29]), .C(C_data_point[29]));
PDUSDGZ I_D_P30 (.PAD(data_point[30]), .C(C_data_point[30]));
PDUSDGZ I_D_P31 (.PAD(data_point[31]), .C(C_data_point[31]));
PDUSDGZ I_D_T0  (.PAD(target[0]),  .C(C_target[0]));
PDUSDGZ I_D_T1  (.PAD(target[1]),  .C(C_target[1]));
PDUSDGZ I_D_T2  (.PAD(target[2]),  .C(C_target[2]));
PDUSDGZ I_D_T3  (.PAD(target[3]),  .C(C_target[3]));
PDUSDGZ I_D_T4  (.PAD(target[4]),  .C(C_target[4]));
PDUSDGZ I_D_T5  (.PAD(target[5]),  .C(C_target[5]));
PDUSDGZ I_D_T6  (.PAD(target[6]),  .C(C_target[6]));
PDUSDGZ I_D_T7  (.PAD(target[7]),  .C(C_target[7]));
PDUSDGZ I_D_T8  (.PAD(target[8]),  .C(C_target[8]));
PDUSDGZ I_D_T9  (.PAD(target[9]),  .C(C_target[9]));
PDUSDGZ I_D_T10 (.PAD(target[10]), .C(C_target[10]));
PDUSDGZ I_D_T11 (.PAD(target[11]), .C(C_target[11]));
PDUSDGZ I_D_T12 (.PAD(target[12]), .C(C_target[12]));
PDUSDGZ I_D_T13 (.PAD(target[13]), .C(C_target[13]));
PDUSDGZ I_D_T14 (.PAD(target[14]), .C(C_target[14]));
PDUSDGZ I_D_T15 (.PAD(target[15]), .C(C_target[15]));
PDUSDGZ I_D_T16 (.PAD(target[16]), .C(C_target[16]));
PDUSDGZ I_D_T17 (.PAD(target[17]), .C(C_target[17]));
PDUSDGZ I_D_T18 (.PAD(target[18]), .C(C_target[18]));
PDUSDGZ I_D_T19 (.PAD(target[19]), .C(C_target[19]));
PDUSDGZ I_D_T20 (.PAD(target[20]), .C(C_target[20]));
PDUSDGZ I_D_T21 (.PAD(target[21]), .C(C_target[21]));
PDUSDGZ I_D_T22 (.PAD(target[22]), .C(C_target[22]));
PDUSDGZ I_D_T23 (.PAD(target[23]), .C(C_target[23]));
PDUSDGZ I_D_T24 (.PAD(target[24]), .C(C_target[24]));
PDUSDGZ I_D_T25 (.PAD(target[25]), .C(C_target[25]));
PDUSDGZ I_D_T26 (.PAD(target[26]), .C(C_target[26]));
PDUSDGZ I_D_T27 (.PAD(target[27]), .C(C_target[27]));
PDUSDGZ I_D_T28 (.PAD(target[28]), .C(C_target[28]));
PDUSDGZ I_D_T29 (.PAD(target[29]), .C(C_target[29]));
PDUSDGZ I_D_T30 (.PAD(target[30]), .C(C_target[30]));
PDUSDGZ I_D_T31 (.PAD(target[31]), .C(C_target[31]));
PDUSDGZ I_D_W10  (.PAD(weight1[0]),  .C(C_weight1[0]));
PDUSDGZ I_D_W11  (.PAD(weight1[1]),  .C(C_weight1[1]));
PDUSDGZ I_D_W12  (.PAD(weight1[2]),  .C(C_weight1[2]));
PDUSDGZ I_D_W13  (.PAD(weight1[3]),  .C(C_weight1[3]));
PDUSDGZ I_D_W14  (.PAD(weight1[4]),  .C(C_weight1[4]));
PDUSDGZ I_D_W15  (.PAD(weight1[5]),  .C(C_weight1[5]));
PDUSDGZ I_D_W16  (.PAD(weight1[6]),  .C(C_weight1[6]));
PDUSDGZ I_D_W17  (.PAD(weight1[7]),  .C(C_weight1[7]));
PDUSDGZ I_D_W18  (.PAD(weight1[8]),  .C(C_weight1[8]));
PDUSDGZ I_D_W19  (.PAD(weight1[9]),  .C(C_weight1[9]));
PDUSDGZ I_D_W110 (.PAD(weight1[10]), .C(C_weight1[10]));
PDUSDGZ I_D_W111 (.PAD(weight1[11]), .C(C_weight1[11]));
PDUSDGZ I_D_W112 (.PAD(weight1[12]), .C(C_weight1[12]));
PDUSDGZ I_D_W113 (.PAD(weight1[13]), .C(C_weight1[13]));
PDUSDGZ I_D_W114 (.PAD(weight1[14]), .C(C_weight1[14]));
PDUSDGZ I_D_W115 (.PAD(weight1[15]), .C(C_weight1[15]));
PDUSDGZ I_D_W116 (.PAD(weight1[16]), .C(C_weight1[16]));
PDUSDGZ I_D_W117 (.PAD(weight1[17]), .C(C_weight1[17]));
PDUSDGZ I_D_W118 (.PAD(weight1[18]), .C(C_weight1[18]));
PDUSDGZ I_D_W119 (.PAD(weight1[19]), .C(C_weight1[19]));
PDUSDGZ I_D_W120 (.PAD(weight1[20]), .C(C_weight1[20]));
PDUSDGZ I_D_W121 (.PAD(weight1[21]), .C(C_weight1[21]));
PDUSDGZ I_D_W122 (.PAD(weight1[22]), .C(C_weight1[22]));
PDUSDGZ I_D_W123 (.PAD(weight1[23]), .C(C_weight1[23]));
PDUSDGZ I_D_W124 (.PAD(weight1[24]), .C(C_weight1[24]));
PDUSDGZ I_D_W125 (.PAD(weight1[25]), .C(C_weight1[25]));
PDUSDGZ I_D_W126 (.PAD(weight1[26]), .C(C_weight1[26]));
PDUSDGZ I_D_W127 (.PAD(weight1[27]), .C(C_weight1[27]));
PDUSDGZ I_D_W128 (.PAD(weight1[28]), .C(C_weight1[28]));
PDUSDGZ I_D_W129 (.PAD(weight1[29]), .C(C_weight1[29]));
PDUSDGZ I_D_W130 (.PAD(weight1[30]), .C(C_weight1[30]));
PDUSDGZ I_D_W131 (.PAD(weight1[31]), .C(C_weight1[31]));
PDUSDGZ I_D_W20  (.PAD(weight2[0]),  .C(C_weight2[0]));
PDUSDGZ I_D_W21  (.PAD(weight2[1]),  .C(C_weight2[1]));
PDUSDGZ I_D_W22  (.PAD(weight2[2]),  .C(C_weight2[2]));
PDUSDGZ I_D_W23  (.PAD(weight2[3]),  .C(C_weight2[3]));
PDUSDGZ I_D_W24  (.PAD(weight2[4]),  .C(C_weight2[4]));
PDUSDGZ I_D_W25  (.PAD(weight2[5]),  .C(C_weight2[5]));
PDUSDGZ I_D_W26  (.PAD(weight2[6]),  .C(C_weight2[6]));
PDUSDGZ I_D_W27  (.PAD(weight2[7]),  .C(C_weight2[7]));
PDUSDGZ I_D_W28  (.PAD(weight2[8]),  .C(C_weight2[8]));
PDUSDGZ I_D_W29  (.PAD(weight2[9]),  .C(C_weight2[9]));
PDUSDGZ I_D_W210 (.PAD(weight2[10]), .C(C_weight2[10]));
PDUSDGZ I_D_W211 (.PAD(weight2[11]), .C(C_weight2[11]));
PDUSDGZ I_D_W212 (.PAD(weight2[12]), .C(C_weight2[12]));
PDUSDGZ I_D_W213 (.PAD(weight2[13]), .C(C_weight2[13]));
PDUSDGZ I_D_W214 (.PAD(weight2[14]), .C(C_weight2[14]));
PDUSDGZ I_D_W215 (.PAD(weight2[15]), .C(C_weight2[15]));
PDUSDGZ I_D_W216 (.PAD(weight2[16]), .C(C_weight2[16]));
PDUSDGZ I_D_W217 (.PAD(weight2[17]), .C(C_weight2[17]));
PDUSDGZ I_D_W218 (.PAD(weight2[18]), .C(C_weight2[18]));
PDUSDGZ I_D_W219 (.PAD(weight2[19]), .C(C_weight2[19]));
PDUSDGZ I_D_W220 (.PAD(weight2[20]), .C(C_weight2[20]));
PDUSDGZ I_D_W221 (.PAD(weight2[21]), .C(C_weight2[21]));
PDUSDGZ I_D_W222 (.PAD(weight2[22]), .C(C_weight2[22]));
PDUSDGZ I_D_W223 (.PAD(weight2[23]), .C(C_weight2[23]));
PDUSDGZ I_D_W224 (.PAD(weight2[24]), .C(C_weight2[24]));
PDUSDGZ I_D_W225 (.PAD(weight2[25]), .C(C_weight2[25]));
PDUSDGZ I_D_W226 (.PAD(weight2[26]), .C(C_weight2[26]));
PDUSDGZ I_D_W227 (.PAD(weight2[27]), .C(C_weight2[27]));
PDUSDGZ I_D_W228 (.PAD(weight2[28]), .C(C_weight2[28]));
PDUSDGZ I_D_W229 (.PAD(weight2[29]), .C(C_weight2[29]));
PDUSDGZ I_D_W230 (.PAD(weight2[30]), .C(C_weight2[30]));
PDUSDGZ I_D_W231 (.PAD(weight2[31]), .C(C_weight2[31]));


// Output Pads
PDD08SDGZ O_OUT_VALID(.OEN(1'b0), .I(C_out_valid), .PAD(out_valid), .C());
PDD08SDGZ O_OUT0  (.OEN(1'b0), .I(C_out[0]),  .PAD(out[0]),  .C());
PDD08SDGZ O_OUT1  (.OEN(1'b0), .I(C_out[1]),  .PAD(out[1]),  .C());
PDD08SDGZ O_OUT2  (.OEN(1'b0), .I(C_out[2]),  .PAD(out[2]),  .C());
PDD08SDGZ O_OUT3  (.OEN(1'b0), .I(C_out[3]),  .PAD(out[3]),  .C());
PDD08SDGZ O_OUT4  (.OEN(1'b0), .I(C_out[4]),  .PAD(out[4]),  .C());
PDD08SDGZ O_OUT5  (.OEN(1'b0), .I(C_out[5]),  .PAD(out[5]),  .C());
PDD08SDGZ O_OUT6  (.OEN(1'b0), .I(C_out[6]),  .PAD(out[6]),  .C());
PDD08SDGZ O_OUT7  (.OEN(1'b0), .I(C_out[7]),  .PAD(out[7]),  .C());
PDD08SDGZ O_OUT8  (.OEN(1'b0), .I(C_out[8]),  .PAD(out[8]),  .C());
PDD08SDGZ O_OUT9  (.OEN(1'b0), .I(C_out[9]),  .PAD(out[9]),  .C());
PDD08SDGZ O_OUT10 (.OEN(1'b0), .I(C_out[10]), .PAD(out[10]), .C());
PDD08SDGZ O_OUT11 (.OEN(1'b0), .I(C_out[11]), .PAD(out[11]), .C());
PDD08SDGZ O_OUT12 (.OEN(1'b0), .I(C_out[12]), .PAD(out[12]), .C());
PDD08SDGZ O_OUT13 (.OEN(1'b0), .I(C_out[13]), .PAD(out[13]), .C());
PDD08SDGZ O_OUT14 (.OEN(1'b0), .I(C_out[14]), .PAD(out[14]), .C());
PDD08SDGZ O_OUT15 (.OEN(1'b0), .I(C_out[15]), .PAD(out[15]), .C());
PDD08SDGZ O_OUT16 (.OEN(1'b0), .I(C_out[16]), .PAD(out[16]), .C());
PDD08SDGZ O_OUT17 (.OEN(1'b0), .I(C_out[17]), .PAD(out[17]), .C());
PDD08SDGZ O_OUT18 (.OEN(1'b0), .I(C_out[18]), .PAD(out[18]), .C());
PDD08SDGZ O_OUT19 (.OEN(1'b0), .I(C_out[19]), .PAD(out[19]), .C());
PDD08SDGZ O_OUT20 (.OEN(1'b0), .I(C_out[20]), .PAD(out[20]), .C());
PDD08SDGZ O_OUT21 (.OEN(1'b0), .I(C_out[21]), .PAD(out[21]), .C());
PDD08SDGZ O_OUT22 (.OEN(1'b0), .I(C_out[22]), .PAD(out[22]), .C());
PDD08SDGZ O_OUT23 (.OEN(1'b0), .I(C_out[23]), .PAD(out[23]), .C());
PDD08SDGZ O_OUT24 (.OEN(1'b0), .I(C_out[24]), .PAD(out[24]), .C());
PDD08SDGZ O_OUT25 (.OEN(1'b0), .I(C_out[25]), .PAD(out[25]), .C());
PDD08SDGZ O_OUT26 (.OEN(1'b0), .I(C_out[26]), .PAD(out[26]), .C());
PDD08SDGZ O_OUT27 (.OEN(1'b0), .I(C_out[27]), .PAD(out[27]), .C());
PDD08SDGZ O_OUT28 (.OEN(1'b0), .I(C_out[28]), .PAD(out[28]), .C());
PDD08SDGZ O_OUT29 (.OEN(1'b0), .I(C_out[29]), .PAD(out[29]), .C());
PDD08SDGZ O_OUT30 (.OEN(1'b0), .I(C_out[30]), .PAD(out[30]), .C());
PDD08SDGZ O_OUT31 (.OEN(1'b0), .I(C_out[31]), .PAD(out[31]), .C());



// IO power 
PVDD2DGZ VDDP0 ();
PVSS2DGZ GNDP0 ();
PVDD2DGZ VDDP1 ();
PVSS2DGZ GNDP1 ();
PVDD2DGZ VDDP2 ();
PVSS2DGZ GNDP2 ();
PVDD2DGZ VDDP3 ();
PVSS2DGZ GNDP3 ();
PVDD2DGZ VDDP4 ();
PVSS2DGZ GNDP4 ();
PVDD2DGZ VDDP5 ();
PVSS2DGZ GNDP5 ();
PVDD2DGZ VDDP6 ();
PVSS2DGZ GNDP6 ();
PVDD2DGZ VDDP7 ();
PVSS2DGZ GNDP7 ();


// Core power
PVDD1DGZ VDDC0 ();
PVSS1DGZ GNDC0 ();
PVDD1DGZ VDDC1 ();
PVSS1DGZ GNDC1 ();
PVDD1DGZ VDDC2 ();
PVSS1DGZ GNDC2 ();
PVDD1DGZ VDDC3 ();
PVSS1DGZ GNDC3 ();
PVDD1DGZ VDDC4 ();
PVSS1DGZ GNDC4 ();
PVDD1DGZ VDDC5 ();
PVSS1DGZ GNDC5 ();
PVDD1DGZ VDDC6 ();
PVSS1DGZ GNDC6 ();
PVDD1DGZ VDDC7 ();
PVSS1DGZ GNDC7 ();

endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : O-2018.06-SP1
// Date      : Sun Nov 30 07:59:13 2025
/////////////////////////////////////////////////////////////


module NN ( clk, rst_n, in_valid_d, in_valid_t, in_valid_w1, in_valid_w2, 
        data_point, target, weight1, weight2, out_valid, out );
  input [31:0] data_point;
  input [31:0] target;
  input [31:0] weight1;
  input [31:0] weight2;
  output [31:0] out;
  input clk, rst_n, in_valid_d, in_valid_t, in_valid_w1, in_valid_w2;
  output out_valid;
  wire   N40, N41, N42, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2633, n2634, n2638, n2639, n2641, n2642, n2643, n2644,
         n2646, n2647, n2648, n2649, n2651, M5_b_18_, M5_a_0_, M5_a_2_,
         M5_a_4_, M5_a_6_, M5_a_8_, M5_a_10_, M5_a_12_, M5_a_18_, M5_a_20_,
         M5_a_22_, M4_a_0_, M4_a_1_, M4_a_2_, M4_a_4_, M4_a_5_, M4_a_6_,
         M4_a_7_, M4_a_9_, M4_a_12_, M4_a_13_, M4_a_17_, M4_a_18_, M4_a_19_,
         M4_a_20_, M3_a_0_, M3_a_2_, M3_a_9_, M3_a_10_, M3_a_11_, M3_a_16_,
         M3_a_20_, M3_a_22_, M2_b_0_, M2_b_2_, M2_b_4_, M2_b_6_, M2_b_7_,
         M2_b_8_, M2_b_10_, M2_b_12_, M2_b_13_, M2_b_15_, M2_b_16_, M2_b_17_,
         M2_b_18_, M2_b_19_, M2_a_0_, M2_a_2_, M2_a_3_, M2_a_4_, M2_a_5_,
         M2_a_6_, M2_a_7_, M2_a_8_, M2_a_10_, M2_a_12_, M2_a_14_, M2_a_16_,
         M2_a_17_, M2_a_18_, M2_a_19_, M2_a_22_, M1_b_0_, M1_b_2_, M1_b_3_,
         M1_b_4_, M1_b_6_, M1_b_8_, M1_b_10_, M1_b_11_, M1_b_12_, M1_b_14_,
         M1_b_15_, M1_b_18_, M1_b_19_, M1_b_20_, M1_b_22_, M1_a_0_, M1_a_1_,
         M1_a_2_, M1_a_3_, M1_a_4_, M1_a_5_, M1_a_6_, M1_a_7_, M1_a_8_,
         M1_a_9_, M1_a_10_, M1_a_11_, M1_a_12_, M1_a_13_, M1_a_14_, M1_a_15_,
         M1_a_16_, M1_a_17_, M1_a_19_, M1_a_20_, M1_a_21_, M1_a_22_, M0_b_0_,
         M0_b_1_, M0_b_2_, M0_b_4_, M0_b_5_, M0_b_6_, M0_b_7_, M0_b_8_,
         M0_b_9_, M0_b_10_, M0_b_11_, M0_b_13_, M0_b_15_, M0_b_17_, M0_b_18_,
         M0_b_20_, M0_b_21_, M0_a_0_, M0_a_2_, M0_a_3_, M0_a_4_, M0_a_6_,
         M0_a_7_, M0_a_8_, M0_a_10_, M0_a_12_, M0_a_15_, M0_a_16_, M0_a_18_,
         M0_a_20_, M0_a_22_, M6_mult_x_15_n1207, M6_mult_x_15_n1206,
         M6_mult_x_15_n1205, M6_mult_x_15_n1204, M6_mult_x_15_n1203,
         M6_mult_x_15_n1202, M6_mult_x_15_n1201, M6_mult_x_15_n1200,
         M6_mult_x_15_n1199, M6_mult_x_15_n1198, M6_mult_x_15_n1197,
         M6_mult_x_15_n1196, M6_mult_x_15_n1195, M6_mult_x_15_n1194,
         M6_mult_x_15_n1193, M6_mult_x_15_n1192, M6_mult_x_15_n1191,
         M6_mult_x_15_n1183, M6_mult_x_15_n1182, M6_mult_x_15_n1181,
         M6_mult_x_15_n1180, M6_mult_x_15_n1179, M6_mult_x_15_n1178,
         M6_mult_x_15_n1177, M6_mult_x_15_n1176, M6_mult_x_15_n1175,
         M6_mult_x_15_n1174, M6_mult_x_15_n1173, M6_mult_x_15_n1172,
         M6_mult_x_15_n1171, M6_mult_x_15_n1170, M6_mult_x_15_n1169,
         M6_mult_x_15_n1168, M6_mult_x_15_n1167, M6_mult_x_15_n1166,
         M6_mult_x_15_n1165, M6_mult_x_15_n1164, M6_mult_x_15_n1159,
         M6_mult_x_15_n1158, M6_mult_x_15_n1157, M6_mult_x_15_n1156,
         M6_mult_x_15_n1155, M6_mult_x_15_n1154, M6_mult_x_15_n1153,
         M6_mult_x_15_n1152, M6_mult_x_15_n1151, M6_mult_x_15_n1150,
         M6_mult_x_15_n1149, M6_mult_x_15_n1148, M6_mult_x_15_n1147,
         M6_mult_x_15_n1146, M6_mult_x_15_n1145, M6_mult_x_15_n1144,
         M6_mult_x_15_n1143, M6_mult_x_15_n1142, M6_mult_x_15_n1141,
         M6_mult_x_15_n1140, M6_mult_x_15_n1139, M6_mult_x_15_n1138,
         M6_mult_x_15_n1137, M6_mult_x_15_n1129, M6_mult_x_15_n1128,
         M6_mult_x_15_n1127, M6_mult_x_15_n1126, M6_mult_x_15_n1125,
         M6_mult_x_15_n1124, M6_mult_x_15_n1123, M6_mult_x_15_n1122,
         M6_mult_x_15_n1121, M6_mult_x_15_n1120, M6_mult_x_15_n1119,
         M6_mult_x_15_n1118, M6_mult_x_15_n1117, M6_mult_x_15_n1116,
         M6_mult_x_15_n1115, M6_mult_x_15_n1114, M6_mult_x_15_n1113,
         M6_mult_x_15_n1112, M6_mult_x_15_n1111, M6_mult_x_15_n1110,
         M6_mult_x_15_n1105, M6_mult_x_15_n1104, M6_mult_x_15_n1103,
         M6_mult_x_15_n1102, M6_mult_x_15_n1101, M6_mult_x_15_n1100,
         M6_mult_x_15_n1099, M6_mult_x_15_n1098, M6_mult_x_15_n1097,
         M6_mult_x_15_n1096, M6_mult_x_15_n1095, M6_mult_x_15_n1094,
         M6_mult_x_15_n1093, M6_mult_x_15_n1092, M6_mult_x_15_n1091,
         M6_mult_x_15_n1090, M6_mult_x_15_n1089, M6_mult_x_15_n1088,
         M6_mult_x_15_n1087, M6_mult_x_15_n1086, M6_mult_x_15_n1085,
         M6_mult_x_15_n1084, M6_mult_x_15_n1083, M6_mult_x_15_n1075,
         M6_mult_x_15_n1074, M6_mult_x_15_n1073, M6_mult_x_15_n1072,
         M6_mult_x_15_n1071, M6_mult_x_15_n1070, M6_mult_x_15_n1069,
         M6_mult_x_15_n1068, M6_mult_x_15_n1067, M6_mult_x_15_n1066,
         M6_mult_x_15_n1065, M6_mult_x_15_n1064, M6_mult_x_15_n1063,
         M6_mult_x_15_n1062, M6_mult_x_15_n1061, M6_mult_x_15_n1060,
         M6_mult_x_15_n1059, M6_mult_x_15_n1058, M6_mult_x_15_n1056,
         M6_mult_x_15_n1051, M6_mult_x_15_n1050, M6_mult_x_15_n1049,
         M6_mult_x_15_n1048, M6_mult_x_15_n1047, M6_mult_x_15_n1046,
         M6_mult_x_15_n1045, M6_mult_x_15_n1044, M6_mult_x_15_n1043,
         M6_mult_x_15_n1042, M6_mult_x_15_n1041, M6_mult_x_15_n1040,
         M6_mult_x_15_n1038, M6_mult_x_15_n1037, M6_mult_x_15_n1036,
         M6_mult_x_15_n1035, M6_mult_x_15_n1034, M6_mult_x_15_n1033,
         M6_mult_x_15_n1032, M6_mult_x_15_n1031, M6_mult_x_15_n1030,
         M6_mult_x_15_n1029, M6_mult_x_15_n1020, M6_mult_x_15_n1019,
         M6_mult_x_15_n1018, M6_mult_x_15_n1017, M6_mult_x_15_n1016,
         M6_mult_x_15_n1014, M6_mult_x_15_n1013, M6_mult_x_15_n1012,
         M6_mult_x_15_n1011, M6_mult_x_15_n1010, M6_mult_x_15_n1008,
         M6_mult_x_15_n1007, M6_mult_x_15_n1006, M6_mult_x_15_n1005,
         M6_mult_x_15_n727, M6_mult_x_15_n724, M6_mult_x_15_n722,
         M6_mult_x_15_n721, M6_mult_x_15_n720, M6_mult_x_15_n719,
         M6_mult_x_15_n717, M6_mult_x_15_n716, M6_mult_x_15_n715,
         M6_mult_x_15_n714, M6_mult_x_15_n712, M6_mult_x_15_n711,
         M6_mult_x_15_n710, M6_mult_x_15_n707, M6_mult_x_15_n705,
         M6_mult_x_15_n704, M6_mult_x_15_n703, M6_mult_x_15_n700,
         M6_mult_x_15_n698, M6_mult_x_15_n697, M6_mult_x_15_n696,
         M6_mult_x_15_n694, M6_mult_x_15_n693, M6_mult_x_15_n692,
         M6_mult_x_15_n691, M6_mult_x_15_n690, M6_mult_x_15_n689,
         M6_mult_x_15_n688, M6_mult_x_15_n686, M6_mult_x_15_n685,
         M6_mult_x_15_n684, M6_mult_x_15_n683, M6_mult_x_15_n682,
         M6_mult_x_15_n681, M6_mult_x_15_n680, M6_mult_x_15_n678,
         M6_mult_x_15_n677, M6_mult_x_15_n676, M6_mult_x_15_n675,
         M6_mult_x_15_n674, M6_mult_x_15_n673, M6_mult_x_15_n672,
         M6_mult_x_15_n670, M6_mult_x_15_n669, M6_mult_x_15_n668,
         M6_mult_x_15_n667, M6_mult_x_15_n666, M6_mult_x_15_n665,
         M6_mult_x_15_n662, M6_mult_x_15_n660, M6_mult_x_15_n659,
         M6_mult_x_15_n658, M6_mult_x_15_n657, M6_mult_x_15_n656,
         M6_mult_x_15_n655, M6_mult_x_15_n652, M6_mult_x_15_n650,
         M6_mult_x_15_n649, M6_mult_x_15_n648, M6_mult_x_15_n647,
         M6_mult_x_15_n646, M6_mult_x_15_n645, M6_mult_x_15_n643,
         M6_mult_x_15_n642, M6_mult_x_15_n641, M6_mult_x_15_n640,
         M6_mult_x_15_n639, M6_mult_x_15_n638, M6_mult_x_15_n637,
         M6_mult_x_15_n636, M6_mult_x_15_n635, M6_mult_x_15_n634,
         M6_mult_x_15_n632, M6_mult_x_15_n631, M6_mult_x_15_n630,
         M6_mult_x_15_n629, M6_mult_x_15_n628, M6_mult_x_15_n627,
         M6_mult_x_15_n626, M6_mult_x_15_n625, M6_mult_x_15_n624,
         M6_mult_x_15_n623, M6_mult_x_15_n621, M6_mult_x_15_n620,
         M6_mult_x_15_n619, M6_mult_x_15_n618, M6_mult_x_15_n617,
         M6_mult_x_15_n616, M6_mult_x_15_n615, M6_mult_x_15_n614,
         M6_mult_x_15_n613, M6_mult_x_15_n612, M6_mult_x_15_n610,
         M6_mult_x_15_n609, M6_mult_x_15_n608, M6_mult_x_15_n607,
         M6_mult_x_15_n606, M6_mult_x_15_n605, M6_mult_x_15_n604,
         M6_mult_x_15_n603, M6_mult_x_15_n602, M6_mult_x_15_n601,
         M6_mult_x_15_n599, M6_mult_x_15_n598, M6_mult_x_15_n597,
         M6_mult_x_15_n596, M6_mult_x_15_n595, M6_mult_x_15_n594,
         M6_mult_x_15_n593, M6_mult_x_15_n592, M6_mult_x_15_n591,
         M6_mult_x_15_n590, M6_mult_x_15_n589, M6_mult_x_15_n588,
         M6_mult_x_15_n587, M6_mult_x_15_n586, M6_mult_x_15_n585,
         M6_mult_x_15_n584, M6_mult_x_15_n583, M6_mult_x_15_n582,
         M6_mult_x_15_n581, M6_mult_x_15_n580, M6_mult_x_15_n579,
         M6_mult_x_15_n578, M6_mult_x_15_n577, M6_mult_x_15_n576,
         M6_mult_x_15_n575, M6_mult_x_15_n574, M6_mult_x_15_n573,
         M6_mult_x_15_n572, M6_mult_x_15_n571, M6_mult_x_15_n570,
         M6_mult_x_15_n569, M6_mult_x_15_n568, M6_mult_x_15_n567,
         M6_mult_x_15_n566, M6_mult_x_15_n565, M6_mult_x_15_n564,
         M6_mult_x_15_n563, M6_mult_x_15_n562, M6_mult_x_15_n561,
         M6_mult_x_15_n560, M6_mult_x_15_n559, M6_mult_x_15_n558,
         M6_mult_x_15_n557, M6_mult_x_15_n556, M6_mult_x_15_n555,
         M6_mult_x_15_n554, M6_mult_x_15_n553, M6_mult_x_15_n552,
         M6_mult_x_15_n551, M6_mult_x_15_n550, M6_mult_x_15_n549,
         M6_mult_x_15_n548, M6_mult_x_15_n547, M6_mult_x_15_n546,
         M6_mult_x_15_n545, M6_mult_x_15_n544, M6_mult_x_15_n543,
         M6_mult_x_15_n542, M6_mult_x_15_n541, M6_mult_x_15_n540,
         M6_mult_x_15_n539, M6_mult_x_15_n538, M6_mult_x_15_n537,
         M6_mult_x_15_n536, M6_mult_x_15_n534, M6_mult_x_15_n533,
         M6_mult_x_15_n532, M6_mult_x_15_n531, M6_mult_x_15_n530,
         M6_mult_x_15_n529, M6_mult_x_15_n528, M6_mult_x_15_n527,
         M6_mult_x_15_n526, M6_mult_x_15_n524, M6_mult_x_15_n523,
         M6_mult_x_15_n522, M6_mult_x_15_n521, M6_mult_x_15_n520,
         M6_mult_x_15_n519, M6_mult_x_15_n518, M6_mult_x_15_n517,
         M6_mult_x_15_n516, M6_mult_x_15_n515, M6_mult_x_15_n514,
         M6_mult_x_15_n513, M6_mult_x_15_n512, M6_mult_x_15_n511,
         M6_mult_x_15_n510, M6_mult_x_15_n509, M6_mult_x_15_n508,
         M6_mult_x_15_n507, M6_mult_x_15_n505, M6_mult_x_15_n504,
         M6_mult_x_15_n503, M6_mult_x_15_n502, M6_mult_x_15_n501,
         M6_mult_x_15_n500, M6_mult_x_15_n499, M6_mult_x_15_n498,
         M6_mult_x_15_n496, M6_mult_x_15_n495, M6_mult_x_15_n494,
         M6_mult_x_15_n493, M6_mult_x_15_n492, M6_mult_x_15_n491,
         M6_mult_x_15_n490, M6_mult_x_15_n489, M6_mult_x_15_n488,
         M6_mult_x_15_n487, M6_mult_x_15_n486, M6_mult_x_15_n485,
         M6_mult_x_15_n484, M6_mult_x_15_n483, M6_mult_x_15_n482,
         M6_mult_x_15_n481, M6_mult_x_15_n479, M6_mult_x_15_n478,
         M6_mult_x_15_n477, M6_mult_x_15_n476, M6_mult_x_15_n475,
         M6_mult_x_15_n474, M6_mult_x_15_n472, M6_mult_x_15_n471,
         M6_mult_x_15_n470, M6_mult_x_15_n469, M6_mult_x_15_n468,
         M6_mult_x_15_n467, M6_mult_x_15_n466, M6_mult_x_15_n465,
         M6_mult_x_15_n464, M6_mult_x_15_n463, M6_mult_x_15_n462,
         M6_mult_x_15_n461, M6_mult_x_15_n459, M6_mult_x_15_n458,
         M6_mult_x_15_n457, M6_mult_x_15_n456, M6_mult_x_15_n455,
         M6_mult_x_15_n453, M6_mult_x_15_n452, M6_mult_x_15_n451,
         M6_mult_x_15_n450, M6_mult_x_15_n449, M6_mult_x_15_n448,
         M6_mult_x_15_n447, M6_mult_x_15_n446, M6_mult_x_15_n445,
         M6_mult_x_15_n444, M6_mult_x_15_n442, M6_mult_x_15_n441,
         M6_mult_x_15_n440, M6_mult_x_15_n438, M6_mult_x_15_n437,
         M6_mult_x_15_n436, M6_mult_x_15_n435, M6_mult_x_15_n434,
         M6_mult_x_15_n433, M2_U3_U1_enc_tree_0__2__28_,
         M2_U3_U1_enc_tree_0__2__20_, M2_U3_U1_enc_tree_0__2__12_,
         M2_U3_U1_enc_tree_0__1__30_, M2_U3_U1_enc_tree_0__1__26_,
         M2_U3_U1_enc_tree_0__1__22_, M2_U3_U1_enc_tree_0__1__18_,
         M2_U3_U1_enc_tree_0__1__14_, M2_U3_U1_enc_tree_0__1__10_,
         M2_U3_U1_or2_tree_0__2__24_, M2_U3_U1_or2_tree_0__2__16_,
         M2_U3_U1_or2_tree_0__1__28_, M2_U3_U1_or2_tree_0__1__24_,
         M2_U3_U1_or2_tree_0__1__20_, M2_U3_U1_or2_tree_0__1__16_,
         M2_U3_U1_or2_tree_0__1__12_, M2_U3_U1_or2_tree_1__2__24_,
         M2_U3_U1_or2_tree_1__2__16_, M2_U3_U1_or2_inv_2__24_,
         M2_U3_U1_or2_inv_1__28_, M2_U3_U1_or2_inv_1__24_,
         M2_U3_U1_or2_inv_1__20_, M2_U3_U1_or2_inv_1__12_,
         M2_U3_U1_or2_inv_0__28_, M2_U3_U1_or2_inv_0__24_,
         M2_U3_U1_or2_inv_0__20_, M2_U3_U1_enc_tree_2__4__16_,
         M2_U3_U1_enc_tree_2__3__24_, M2_U3_U1_enc_tree_2__2__28_,
         M2_U3_U1_enc_tree_2__2__24_, M2_U3_U1_enc_tree_2__2__20_,
         M2_U3_U1_enc_tree_2__2__16_, M2_U3_U1_enc_tree_1__4__16_,
         M2_U3_U1_enc_tree_1__3__24_, M2_U3_U1_enc_tree_1__3__8_,
         M2_U3_U1_enc_tree_1__2__28_, M2_U3_U1_enc_tree_1__2__20_,
         M2_U3_U1_enc_tree_1__2__12_, M2_U3_U1_enc_tree_1__1__30_,
         M2_U3_U1_enc_tree_1__1__28_, M2_U3_U1_enc_tree_1__1__26_,
         M2_U3_U1_enc_tree_1__1__24_, M2_U3_U1_enc_tree_1__1__22_,
         M2_U3_U1_enc_tree_1__1__20_, M2_U3_U1_enc_tree_1__1__18_,
         M2_U3_U1_enc_tree_1__1__16_, M2_U3_U1_enc_tree_1__1__14_,
         M2_U3_U1_enc_tree_1__1__12_, M2_U3_U1_enc_tree_1__1__10_,
         M2_U3_U1_enc_tree_0__4__16_, M2_U3_U1_enc_tree_0__3__24_,
         M2_U3_U1_enc_tree_0__3__8_, M2_U3_U1_enc_tree_4__4__16_,
         M2_U3_U1_enc_tree_3__3__24_, M2_U3_U1_enc_tree_3__3__16_,
         M1_U3_U1_enc_tree_0__2__28_, M1_U3_U1_enc_tree_0__2__20_,
         M1_U3_U1_enc_tree_0__2__12_, M1_U3_U1_enc_tree_0__1__30_,
         M1_U3_U1_enc_tree_0__1__26_, M1_U3_U1_enc_tree_0__1__22_,
         M1_U3_U1_enc_tree_0__1__18_, M1_U3_U1_enc_tree_0__1__14_,
         M1_U3_U1_enc_tree_0__1__10_, M1_U3_U1_or2_tree_0__2__24_,
         M1_U3_U1_or2_tree_0__2__16_, M1_U3_U1_or2_tree_0__1__28_,
         M1_U3_U1_or2_tree_0__1__24_, M1_U3_U1_or2_tree_0__1__20_,
         M1_U3_U1_or2_tree_0__1__16_, M1_U3_U1_or2_tree_0__1__12_,
         M1_U3_U1_or2_tree_1__2__24_, M1_U3_U1_or2_tree_1__2__16_,
         M1_U3_U1_or2_inv_2__24_, M1_U3_U1_or2_inv_1__28_,
         M1_U3_U1_or2_inv_1__24_, M1_U3_U1_or2_inv_1__20_,
         M1_U3_U1_or2_inv_1__12_, M1_U3_U1_or2_inv_0__28_,
         M1_U3_U1_or2_inv_0__26_, M1_U3_U1_or2_inv_0__24_,
         M1_U3_U1_or2_inv_0__22_, M1_U3_U1_or2_inv_0__20_,
         M1_U3_U1_or2_inv_0__18_, M1_U3_U1_or2_inv_0__14_,
         M1_U3_U1_or2_inv_0__10_, M1_U3_U1_enc_tree_2__4__16_,
         M1_U3_U1_enc_tree_2__3__24_, M1_U3_U1_enc_tree_2__2__28_,
         M1_U3_U1_enc_tree_2__2__24_, M1_U3_U1_enc_tree_2__2__20_,
         M1_U3_U1_enc_tree_2__2__16_, M1_U3_U1_enc_tree_1__4__16_,
         M1_U3_U1_enc_tree_1__3__24_, M1_U3_U1_enc_tree_1__3__8_,
         M1_U3_U1_enc_tree_1__2__28_, M1_U3_U1_enc_tree_1__2__20_,
         M1_U3_U1_enc_tree_1__2__12_, M1_U3_U1_enc_tree_1__1__30_,
         M1_U3_U1_enc_tree_1__1__28_, M1_U3_U1_enc_tree_1__1__26_,
         M1_U3_U1_enc_tree_1__1__24_, M1_U3_U1_enc_tree_1__1__22_,
         M1_U3_U1_enc_tree_1__1__20_, M1_U3_U1_enc_tree_1__1__18_,
         M1_U3_U1_enc_tree_1__1__16_, M1_U3_U1_enc_tree_1__1__14_,
         M1_U3_U1_enc_tree_1__1__12_, M1_U3_U1_enc_tree_1__1__10_,
         M1_U3_U1_enc_tree_0__4__16_, M1_U3_U1_enc_tree_0__3__24_,
         M1_U3_U1_enc_tree_0__3__8_, M1_U3_U1_enc_tree_3__3__24_,
         M1_U3_U1_enc_tree_3__3__16_, M2_U4_U1_enc_tree_0__2__28_,
         M2_U4_U1_enc_tree_0__2__20_, M2_U4_U1_enc_tree_0__2__12_,
         M2_U4_U1_enc_tree_0__1__30_, M2_U4_U1_enc_tree_0__1__26_,
         M2_U4_U1_enc_tree_0__1__22_, M2_U4_U1_enc_tree_0__1__18_,
         M2_U4_U1_enc_tree_0__1__14_, M2_U4_U1_enc_tree_0__1__10_,
         M2_U4_U1_or2_tree_0__2__24_, M2_U4_U1_or2_tree_0__2__16_,
         M2_U4_U1_or2_tree_0__1__28_, M2_U4_U1_or2_tree_0__1__24_,
         M2_U4_U1_or2_tree_0__1__20_, M2_U4_U1_or2_tree_0__1__16_,
         M2_U4_U1_or2_tree_1__2__24_, M2_U4_U1_or2_tree_1__2__16_,
         M2_U4_U1_or2_inv_2__24_, M2_U4_U1_or2_inv_1__28_,
         M2_U4_U1_or2_inv_1__24_, M2_U4_U1_or2_inv_1__20_,
         M2_U4_U1_or2_inv_1__12_, M2_U4_U1_or2_inv_0__28_,
         M2_U4_U1_or2_inv_0__26_, M2_U4_U1_or2_inv_0__24_,
         M2_U4_U1_or2_inv_0__22_, M2_U4_U1_or2_inv_0__20_,
         M2_U4_U1_or2_inv_0__18_, M2_U4_U1_or2_inv_0__14_,
         M2_U4_U1_or2_inv_0__10_, M2_U4_U1_enc_tree_2__4__16_,
         M2_U4_U1_enc_tree_2__3__24_, M2_U4_U1_enc_tree_2__2__28_,
         M2_U4_U1_enc_tree_2__2__24_, M2_U4_U1_enc_tree_2__2__20_,
         M2_U4_U1_enc_tree_2__2__16_, M2_U4_U1_enc_tree_1__4__16_,
         M2_U4_U1_enc_tree_1__3__24_, M2_U4_U1_enc_tree_1__3__8_,
         M2_U4_U1_enc_tree_1__2__28_, M2_U4_U1_enc_tree_1__2__20_,
         M2_U4_U1_enc_tree_1__2__12_, M2_U4_U1_enc_tree_1__1__30_,
         M2_U4_U1_enc_tree_1__1__28_, M2_U4_U1_enc_tree_1__1__26_,
         M2_U4_U1_enc_tree_1__1__24_, M2_U4_U1_enc_tree_1__1__22_,
         M2_U4_U1_enc_tree_1__1__20_, M2_U4_U1_enc_tree_1__1__18_,
         M2_U4_U1_enc_tree_1__1__16_, M2_U4_U1_enc_tree_1__1__14_,
         M2_U4_U1_enc_tree_1__1__12_, M2_U4_U1_enc_tree_1__1__10_,
         M2_U4_U1_enc_tree_0__4__16_, M2_U4_U1_enc_tree_0__3__24_,
         M2_U4_U1_enc_tree_0__3__8_, M2_U4_U1_enc_tree_3__3__24_,
         M2_U4_U1_enc_tree_3__3__16_, M0_U4_U1_enc_tree_0__2__28_,
         M0_U4_U1_enc_tree_0__2__20_, M0_U4_U1_enc_tree_0__2__12_,
         M0_U4_U1_enc_tree_0__1__30_, M0_U4_U1_enc_tree_0__1__26_,
         M0_U4_U1_enc_tree_0__1__22_, M0_U4_U1_enc_tree_0__1__18_,
         M0_U4_U1_enc_tree_0__1__14_, M0_U4_U1_enc_tree_0__1__10_,
         M0_U4_U1_or2_tree_0__2__24_, M0_U4_U1_or2_tree_0__2__16_,
         M0_U4_U1_or2_tree_0__1__28_, M0_U4_U1_or2_tree_0__1__24_,
         M0_U4_U1_or2_tree_0__1__20_, M0_U4_U1_or2_tree_0__1__16_,
         M0_U4_U1_or2_tree_0__1__12_, M0_U4_U1_or2_tree_1__2__24_,
         M0_U4_U1_or2_tree_1__2__16_, M0_U4_U1_or2_inv_2__24_,
         M0_U4_U1_or2_inv_1__24_, M0_U4_U1_or2_inv_1__20_,
         M0_U4_U1_or2_inv_1__12_, M0_U4_U1_or2_inv_0__26_,
         M0_U4_U1_or2_inv_0__24_, M0_U4_U1_or2_inv_0__22_,
         M0_U4_U1_or2_inv_0__20_, M0_U4_U1_or2_inv_0__18_,
         M0_U4_U1_or2_inv_0__14_, M0_U4_U1_or2_inv_0__10_,
         M0_U4_U1_enc_tree_2__4__16_, M0_U4_U1_enc_tree_2__3__24_,
         M0_U4_U1_enc_tree_2__2__28_, M0_U4_U1_enc_tree_2__2__24_,
         M0_U4_U1_enc_tree_2__2__20_, M0_U4_U1_enc_tree_2__2__16_,
         M0_U4_U1_enc_tree_1__4__16_, M0_U4_U1_enc_tree_1__3__24_,
         M0_U4_U1_enc_tree_1__3__8_, M0_U4_U1_enc_tree_1__2__28_,
         M0_U4_U1_enc_tree_1__2__20_, M0_U4_U1_enc_tree_1__2__12_,
         M0_U4_U1_enc_tree_1__1__30_, M0_U4_U1_enc_tree_1__1__28_,
         M0_U4_U1_enc_tree_1__1__26_, M0_U4_U1_enc_tree_1__1__24_,
         M0_U4_U1_enc_tree_1__1__22_, M0_U4_U1_enc_tree_1__1__20_,
         M0_U4_U1_enc_tree_1__1__18_, M0_U4_U1_enc_tree_1__1__16_,
         M0_U4_U1_enc_tree_1__1__14_, M0_U4_U1_enc_tree_1__1__12_,
         M0_U4_U1_enc_tree_1__1__10_, M0_U4_U1_enc_tree_0__4__16_,
         M0_U4_U1_enc_tree_0__3__24_, M0_U4_U1_enc_tree_0__3__8_,
         M0_U4_U1_enc_tree_3__3__24_, M0_U4_U1_enc_tree_3__3__16_,
         M1_U4_U1_enc_tree_0__2__28_, M1_U4_U1_enc_tree_0__2__20_,
         M1_U4_U1_enc_tree_0__2__12_, M1_U4_U1_enc_tree_0__1__30_,
         M1_U4_U1_enc_tree_0__1__26_, M1_U4_U1_enc_tree_0__1__22_,
         M1_U4_U1_enc_tree_0__1__18_, M1_U4_U1_enc_tree_0__1__14_,
         M1_U4_U1_enc_tree_0__1__10_, M1_U4_U1_or2_tree_0__2__24_,
         M1_U4_U1_or2_tree_0__2__16_, M1_U4_U1_or2_tree_0__1__28_,
         M1_U4_U1_or2_tree_0__1__24_, M1_U4_U1_or2_tree_0__1__20_,
         M1_U4_U1_or2_tree_0__1__16_, M1_U4_U1_or2_tree_0__1__12_,
         M1_U4_U1_or2_tree_1__2__24_, M1_U4_U1_or2_tree_1__2__16_,
         M1_U4_U1_or2_inv_2__24_, M1_U4_U1_or2_inv_1__28_,
         M1_U4_U1_or2_inv_1__24_, M1_U4_U1_or2_inv_1__20_,
         M1_U4_U1_or2_inv_1__12_, M1_U4_U1_or2_inv_0__28_,
         M1_U4_U1_or2_inv_0__24_, M1_U4_U1_or2_inv_0__20_,
         M1_U4_U1_enc_tree_2__4__16_, M1_U4_U1_enc_tree_2__3__24_,
         M1_U4_U1_enc_tree_2__2__28_, M1_U4_U1_enc_tree_2__2__24_,
         M1_U4_U1_enc_tree_2__2__20_, M1_U4_U1_enc_tree_2__2__16_,
         M1_U4_U1_enc_tree_1__4__16_, M1_U4_U1_enc_tree_1__3__24_,
         M1_U4_U1_enc_tree_1__3__8_, M1_U4_U1_enc_tree_1__2__28_,
         M1_U4_U1_enc_tree_1__2__20_, M1_U4_U1_enc_tree_1__2__12_,
         M1_U4_U1_enc_tree_1__1__30_, M1_U4_U1_enc_tree_1__1__28_,
         M1_U4_U1_enc_tree_1__1__26_, M1_U4_U1_enc_tree_1__1__24_,
         M1_U4_U1_enc_tree_1__1__22_, M1_U4_U1_enc_tree_1__1__20_,
         M1_U4_U1_enc_tree_1__1__18_, M1_U4_U1_enc_tree_1__1__16_,
         M1_U4_U1_enc_tree_1__1__14_, M1_U4_U1_enc_tree_1__1__12_,
         M1_U4_U1_enc_tree_1__1__10_, M1_U4_U1_enc_tree_0__4__16_,
         M1_U4_U1_enc_tree_0__3__24_, M1_U4_U1_enc_tree_0__3__8_,
         M1_U4_U1_enc_tree_3__3__24_, M1_U4_U1_enc_tree_3__3__16_,
         M0_U3_U1_enc_tree_0__2__28_, M0_U3_U1_enc_tree_0__2__20_,
         M0_U3_U1_enc_tree_0__2__12_, M0_U3_U1_enc_tree_0__1__30_,
         M0_U3_U1_enc_tree_0__1__26_, M0_U3_U1_enc_tree_0__1__22_,
         M0_U3_U1_enc_tree_0__1__18_, M0_U3_U1_enc_tree_0__1__14_,
         M0_U3_U1_enc_tree_0__1__10_, M0_U3_U1_or2_tree_0__2__24_,
         M0_U3_U1_or2_tree_0__2__16_, M0_U3_U1_or2_tree_0__1__28_,
         M0_U3_U1_or2_tree_0__1__24_, M0_U3_U1_or2_tree_0__1__20_,
         M0_U3_U1_or2_tree_0__1__16_, M0_U3_U1_or2_tree_0__1__12_,
         M0_U3_U1_or2_tree_1__2__24_, M0_U3_U1_or2_tree_1__2__16_,
         M0_U3_U1_or2_inv_2__24_, M0_U3_U1_or2_inv_1__28_,
         M0_U3_U1_or2_inv_1__24_, M0_U3_U1_or2_inv_1__20_,
         M0_U3_U1_or2_inv_1__12_, M0_U3_U1_or2_inv_0__28_,
         M0_U3_U1_or2_inv_0__24_, M0_U3_U1_or2_inv_0__20_,
         M0_U3_U1_enc_tree_2__4__16_, M0_U3_U1_enc_tree_2__3__24_,
         M0_U3_U1_enc_tree_2__2__28_, M0_U3_U1_enc_tree_2__2__24_,
         M0_U3_U1_enc_tree_2__2__20_, M0_U3_U1_enc_tree_2__2__16_,
         M0_U3_U1_enc_tree_1__4__16_, M0_U3_U1_enc_tree_1__3__24_,
         M0_U3_U1_enc_tree_1__3__8_, M0_U3_U1_enc_tree_1__2__28_,
         M0_U3_U1_enc_tree_1__2__20_, M0_U3_U1_enc_tree_1__2__12_,
         M0_U3_U1_enc_tree_1__1__30_, M0_U3_U1_enc_tree_1__1__28_,
         M0_U3_U1_enc_tree_1__1__26_, M0_U3_U1_enc_tree_1__1__24_,
         M0_U3_U1_enc_tree_1__1__22_, M0_U3_U1_enc_tree_1__1__20_,
         M0_U3_U1_enc_tree_1__1__18_, M0_U3_U1_enc_tree_1__1__16_,
         M0_U3_U1_enc_tree_1__1__14_, M0_U3_U1_enc_tree_1__1__12_,
         M0_U3_U1_enc_tree_1__1__10_, M0_U3_U1_enc_tree_0__4__16_,
         M0_U3_U1_enc_tree_0__3__24_, M0_U3_U1_enc_tree_0__3__8_,
         M0_U3_U1_enc_tree_3__3__24_, M0_U3_U1_enc_tree_3__3__16_,
         M4_U3_U1_enc_tree_0__2__28_, M4_U3_U1_enc_tree_0__2__20_,
         M4_U3_U1_enc_tree_0__2__12_, M4_U3_U1_enc_tree_0__1__30_,
         M4_U3_U1_enc_tree_0__1__26_, M4_U3_U1_enc_tree_0__1__22_,
         M4_U3_U1_enc_tree_0__1__18_, M4_U3_U1_enc_tree_0__1__14_,
         M4_U3_U1_enc_tree_0__1__10_, M4_U3_U1_or2_tree_0__2__24_,
         M4_U3_U1_or2_tree_0__2__16_, M4_U3_U1_or2_tree_0__1__28_,
         M4_U3_U1_or2_tree_0__1__24_, M4_U3_U1_or2_tree_0__1__20_,
         M4_U3_U1_or2_tree_0__1__16_, M4_U3_U1_or2_tree_0__1__12_,
         M4_U3_U1_or2_tree_1__2__24_, M4_U3_U1_or2_tree_1__2__16_,
         M4_U3_U1_or2_inv_2__24_, M4_U3_U1_or2_inv_1__28_,
         M4_U3_U1_or2_inv_1__24_, M4_U3_U1_or2_inv_1__20_,
         M4_U3_U1_or2_inv_1__12_, M4_U3_U1_or2_inv_0__30_,
         M4_U3_U1_or2_inv_0__28_, M4_U3_U1_or2_inv_0__24_,
         M4_U3_U1_or2_inv_0__20_, M4_U3_U1_enc_tree_2__4__16_,
         M4_U3_U1_enc_tree_2__3__24_, M4_U3_U1_enc_tree_2__2__28_,
         M4_U3_U1_enc_tree_2__2__24_, M4_U3_U1_enc_tree_2__2__20_,
         M4_U3_U1_enc_tree_2__2__16_, M4_U3_U1_enc_tree_1__4__16_,
         M4_U3_U1_enc_tree_1__3__24_, M4_U3_U1_enc_tree_1__3__8_,
         M4_U3_U1_enc_tree_1__2__28_, M4_U3_U1_enc_tree_1__2__20_,
         M4_U3_U1_enc_tree_1__2__12_, M4_U3_U1_enc_tree_1__1__30_,
         M4_U3_U1_enc_tree_1__1__28_, M4_U3_U1_enc_tree_1__1__26_,
         M4_U3_U1_enc_tree_1__1__24_, M4_U3_U1_enc_tree_1__1__22_,
         M4_U3_U1_enc_tree_1__1__20_, M4_U3_U1_enc_tree_1__1__18_,
         M4_U3_U1_enc_tree_1__1__16_, M4_U3_U1_enc_tree_1__1__14_,
         M4_U3_U1_enc_tree_1__1__12_, M4_U3_U1_enc_tree_1__1__10_,
         M4_U3_U1_enc_tree_0__4__16_, M4_U3_U1_enc_tree_0__3__24_,
         M4_U3_U1_enc_tree_0__3__8_, M4_U3_U1_enc_tree_3__3__24_,
         M4_U3_U1_enc_tree_3__3__16_, M3_U3_U1_enc_tree_0__2__28_,
         M3_U3_U1_enc_tree_0__2__20_, M3_U3_U1_enc_tree_0__2__12_,
         M3_U3_U1_enc_tree_0__1__30_, M3_U3_U1_enc_tree_0__1__26_,
         M3_U3_U1_enc_tree_0__1__22_, M3_U3_U1_enc_tree_0__1__18_,
         M3_U3_U1_enc_tree_0__1__14_, M3_U3_U1_enc_tree_0__1__10_,
         M3_U3_U1_or2_tree_0__2__24_, M3_U3_U1_or2_tree_0__2__16_,
         M3_U3_U1_or2_tree_0__1__28_, M3_U3_U1_or2_tree_0__1__24_,
         M3_U3_U1_or2_tree_0__1__20_, M3_U3_U1_or2_tree_0__1__16_,
         M3_U3_U1_or2_tree_1__2__24_, M3_U3_U1_or2_tree_1__2__16_,
         M3_U3_U1_or2_inv_2__24_, M3_U3_U1_or2_inv_1__28_,
         M3_U3_U1_or2_inv_1__24_, M3_U3_U1_or2_inv_1__20_,
         M3_U3_U1_or2_inv_1__12_, M3_U3_U1_or2_inv_0__28_,
         M3_U3_U1_or2_inv_0__24_, M3_U3_U1_or2_inv_0__20_,
         M3_U3_U1_or2_inv_0__18_, M3_U3_U1_enc_tree_2__4__16_,
         M3_U3_U1_enc_tree_2__3__24_, M3_U3_U1_enc_tree_2__2__28_,
         M3_U3_U1_enc_tree_2__2__24_, M3_U3_U1_enc_tree_2__2__20_,
         M3_U3_U1_enc_tree_2__2__16_, M3_U3_U1_enc_tree_1__4__16_,
         M3_U3_U1_enc_tree_1__3__24_, M3_U3_U1_enc_tree_1__3__8_,
         M3_U3_U1_enc_tree_1__2__28_, M3_U3_U1_enc_tree_1__2__20_,
         M3_U3_U1_enc_tree_1__2__12_, M3_U3_U1_enc_tree_1__1__30_,
         M3_U3_U1_enc_tree_1__1__28_, M3_U3_U1_enc_tree_1__1__26_,
         M3_U3_U1_enc_tree_1__1__24_, M3_U3_U1_enc_tree_1__1__22_,
         M3_U3_U1_enc_tree_1__1__20_, M3_U3_U1_enc_tree_1__1__18_,
         M3_U3_U1_enc_tree_1__1__16_, M3_U3_U1_enc_tree_1__1__14_,
         M3_U3_U1_enc_tree_1__1__12_, M3_U3_U1_enc_tree_1__1__10_,
         M3_U3_U1_enc_tree_0__4__16_, M3_U3_U1_enc_tree_0__3__24_,
         M3_U3_U1_enc_tree_0__3__8_, M3_U3_U1_enc_tree_3__3__24_,
         M3_U3_U1_enc_tree_3__3__16_, M5_U3_U1_enc_tree_0__2__28_,
         M5_U3_U1_enc_tree_0__2__20_, M5_U3_U1_enc_tree_0__2__12_,
         M5_U3_U1_enc_tree_0__1__30_, M5_U3_U1_enc_tree_0__1__26_,
         M5_U3_U1_enc_tree_0__1__22_, M5_U3_U1_enc_tree_0__1__18_,
         M5_U3_U1_enc_tree_0__1__14_, M5_U3_U1_enc_tree_0__1__10_,
         M5_U3_U1_or2_tree_0__2__24_, M5_U3_U1_or2_tree_0__2__16_,
         M5_U3_U1_or2_tree_0__1__28_, M5_U3_U1_or2_tree_0__1__24_,
         M5_U3_U1_or2_tree_0__1__20_, M5_U3_U1_or2_tree_0__1__16_,
         M5_U3_U1_or2_tree_1__2__24_, M5_U3_U1_or2_tree_1__2__16_,
         M5_U3_U1_or2_inv_2__24_, M5_U3_U1_or2_inv_1__28_,
         M5_U3_U1_or2_inv_1__24_, M5_U3_U1_or2_inv_1__20_,
         M5_U3_U1_or2_inv_1__12_, M5_U3_U1_or2_inv_0__28_,
         M5_U3_U1_or2_inv_0__24_, M5_U3_U1_or2_inv_0__20_,
         M5_U3_U1_enc_tree_2__4__16_, M5_U3_U1_enc_tree_2__3__24_,
         M5_U3_U1_enc_tree_2__2__28_, M5_U3_U1_enc_tree_2__2__24_,
         M5_U3_U1_enc_tree_2__2__20_, M5_U3_U1_enc_tree_2__2__16_,
         M5_U3_U1_enc_tree_1__4__16_, M5_U3_U1_enc_tree_1__3__24_,
         M5_U3_U1_enc_tree_1__3__8_, M5_U3_U1_enc_tree_1__2__28_,
         M5_U3_U1_enc_tree_1__2__20_, M5_U3_U1_enc_tree_1__2__12_,
         M5_U3_U1_enc_tree_1__1__30_, M5_U3_U1_enc_tree_1__1__28_,
         M5_U3_U1_enc_tree_1__1__26_, M5_U3_U1_enc_tree_1__1__24_,
         M5_U3_U1_enc_tree_1__1__22_, M5_U3_U1_enc_tree_1__1__20_,
         M5_U3_U1_enc_tree_1__1__18_, M5_U3_U1_enc_tree_1__1__16_,
         M5_U3_U1_enc_tree_1__1__14_, M5_U3_U1_enc_tree_1__1__12_,
         M5_U3_U1_enc_tree_1__1__10_, M5_U3_U1_enc_tree_0__4__16_,
         M5_U3_U1_enc_tree_0__3__24_, M5_U3_U1_enc_tree_0__3__8_,
         M5_U3_U1_enc_tree_3__3__24_, M5_U3_U1_enc_tree_3__3__16_,
         M4_U4_U1_enc_tree_0__2__12_, M4_U4_U1_enc_tree_0__1__14_,
         M4_U4_U1_enc_tree_0__1__10_, M4_U4_U1_or2_tree_0__1__28_,
         M4_U4_U1_or2_tree_0__1__24_, M4_U4_U1_or2_tree_0__1__20_,
         M4_U4_U1_or2_tree_0__1__16_, M4_U4_U1_or2_tree_0__1__12_,
         M4_U4_U1_or2_inv_1__12_, M4_U4_U1_or2_inv_0__14_,
         M4_U4_U1_or2_inv_0__10_, M4_U4_U1_enc_tree_2__2__28_,
         M4_U4_U1_enc_tree_2__2__24_, M4_U4_U1_enc_tree_2__2__20_,
         M4_U4_U1_enc_tree_2__2__16_, M4_U4_U1_enc_tree_1__2__12_,
         M4_U4_U1_enc_tree_1__1__30_, M4_U4_U1_enc_tree_1__1__28_,
         M4_U4_U1_enc_tree_1__1__26_, M4_U4_U1_enc_tree_1__1__24_,
         M4_U4_U1_enc_tree_1__1__22_, M4_U4_U1_enc_tree_1__1__20_,
         M4_U4_U1_enc_tree_1__1__18_, M4_U4_U1_enc_tree_1__1__16_,
         M4_U4_U1_enc_tree_1__1__14_, M4_U4_U1_enc_tree_1__1__12_,
         M4_U4_U1_enc_tree_1__1__10_, M4_U4_U1_enc_tree_3__3__24_,
         M4_U4_U1_enc_tree_3__3__16_, M3_U4_U1_enc_tree_0__2__28_,
         M3_U4_U1_enc_tree_0__2__20_, M3_U4_U1_enc_tree_0__1__30_,
         M3_U4_U1_enc_tree_0__1__26_, M3_U4_U1_enc_tree_0__1__22_,
         M3_U4_U1_enc_tree_0__1__18_, M3_U4_U1_or2_tree_0__2__24_,
         M3_U4_U1_or2_tree_0__2__16_, M3_U4_U1_or2_tree_1__2__24_,
         M3_U4_U1_or2_tree_1__2__16_, M3_U4_U1_or2_inv_2__24_,
         M3_U4_U1_or2_inv_1__28_, M3_U4_U1_or2_inv_1__24_,
         M3_U4_U1_or2_inv_1__20_, M3_U4_U1_or2_inv_0__28_,
         M3_U4_U1_or2_inv_0__24_, M3_U4_U1_or2_inv_0__20_,
         M3_U4_U1_or2_inv_0__18_, M3_U4_U1_enc_tree_2__4__16_,
         M3_U4_U1_enc_tree_2__3__24_, M3_U4_U1_enc_tree_1__4__16_,
         M3_U4_U1_enc_tree_1__3__24_, M3_U4_U1_enc_tree_1__3__8_,
         M3_U4_U1_enc_tree_1__2__28_, M3_U4_U1_enc_tree_1__2__20_,
         M3_U4_U1_enc_tree_0__4__16_, M3_U4_U1_enc_tree_0__3__24_,
         M3_U4_U1_enc_tree_0__3__8_, M2_mult_x_15_a_1_, M2_mult_x_15_n1669,
         M2_mult_x_15_n1668, M2_mult_x_15_n43, M3_mult_x_15_b_22_,
         M3_mult_x_15_b_21_, M3_mult_x_15_b_20_, M3_mult_x_15_b_19_,
         M3_mult_x_15_b_17_, M3_mult_x_15_b_15_, M3_mult_x_15_b_14_,
         M3_mult_x_15_b_13_, M3_mult_x_15_b_12_, M3_mult_x_15_b_11_,
         M3_mult_x_15_b_9_, M3_mult_x_15_b_7_, M3_mult_x_15_b_6_,
         M3_mult_x_15_b_5_, M3_mult_x_15_b_3_, M3_mult_x_15_b_2_,
         M3_mult_x_15_b_1_, M3_mult_x_15_a_1_, M3_mult_x_15_a_15_,
         M3_mult_x_15_a_17_, M3_mult_x_15_n1682, M3_mult_x_15_n61,
         M5_mult_x_15_n1, M4_mult_x_15_n1680, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25935, n25936, n25937, n25938, n25939, n25940,
         n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948,
         n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956,
         n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
         n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972,
         n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980,
         n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988,
         n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996,
         n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004,
         n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012,
         n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020,
         n26021, n26024, n26025, n26026, n26027, n26030, n26031, n26032,
         n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
         n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,
         n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
         n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064,
         n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
         n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
         n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088,
         n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
         n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
         n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
         n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
         n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
         n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
         n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,
         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
         n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
         n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,
         n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
         n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
         n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
         n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
         n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
         n26234, n26235, n26239, n26240, n26242, n26243, n26244, n26245,
         n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253,
         n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
         n26262, n26264, n26265, n26266, n26267, n26269, n26270, n26271,
         n26272, n26273, n26274, n26275, n26276, n26277, n26279, n26280,
         n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
         n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,
         n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304,
         n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
         n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
         n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,
         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,
         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,
         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
         n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,
         n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,
         n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
         n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
         n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
         n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
         n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,
         n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
         n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,
         n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520,
         n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528,
         n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,
         n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544,
         n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
         n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
         n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,
         n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
         n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584,
         n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,
         n26593, n26594, n26595;
  wire   [31:0] mul5_out;
  wire   [30:0] learning_rate;
  wire   [31:0] y10;
  wire   [31:0] y11;
  wire   [2:0] cs;
  wire   [2:0] valid;
  wire   [31:0] y12;
  wire   [31:0] temp0;
  wire   [31:0] temp1;
  wire   [31:0] temp2;
  wire   [31:0] y20;
  wire   [31:0] sigma11;
  wire   [31:0] sigma12;
  wire   [31:9] sigma10;
  wire   [31:0] target_temp;
  wire   [95:0] w2;
  wire   [383:0] w1;
  wire   [31:0] temp3;
  wire   [127:0] data;
  wire   [8:0] iter;

  DFFHQXL temp0_reg_30_ ( .D(n2556), .CK(clk), .Q(temp0[30]) );
  DFFHQXL temp0_reg_25_ ( .D(n2566), .CK(clk), .Q(temp0[25]) );
  DFFHQXL temp0_reg_23_ ( .D(n2570), .CK(clk), .Q(temp0[23]) );
  DFFHQXL temp3_reg_30_ ( .D(mul5_out[30]), .CK(clk), .Q(temp3[30]) );
  DFFHQXL temp3_reg_29_ ( .D(mul5_out[29]), .CK(clk), .Q(temp3[29]) );
  DFFHQXL temp3_reg_28_ ( .D(mul5_out[28]), .CK(clk), .Q(temp3[28]) );
  DFFHQXL temp3_reg_27_ ( .D(mul5_out[27]), .CK(clk), .Q(temp3[27]) );
  DFFHQXL temp3_reg_26_ ( .D(mul5_out[26]), .CK(clk), .Q(temp3[26]) );
  DFFHQXL temp3_reg_25_ ( .D(mul5_out[25]), .CK(clk), .Q(temp3[25]) );
  DFFHQXL temp3_reg_23_ ( .D(mul5_out[23]), .CK(clk), .Q(temp3[23]) );
  DFFSX4 cs_reg_0_ ( .D(n2491), .CK(clk), .SN(rst_n), .Q(n26140), .QN(cs[0])
         );
  DFFSX4 cs_reg_1_ ( .D(n2490), .CK(clk), .SN(rst_n), .Q(n25887), .QN(cs[1])
         );
  DFFSX1 y20_reg_31_ ( .D(n2391), .CK(clk), .SN(rst_n), .QN(y20[31]) );
  DFFSX1 target_temp_reg_30_ ( .D(n2262), .CK(clk), .SN(rst_n), .Q(n6173), 
        .QN(target_temp[30]) );
  DFFSX1 target_temp_reg_28_ ( .D(n2260), .CK(clk), .SN(rst_n), .Q(n6170), 
        .QN(target_temp[28]) );
  DFFSX1 target_temp_reg_27_ ( .D(n2259), .CK(clk), .SN(rst_n), .Q(n6171), 
        .QN(target_temp[27]) );
  DFFSX1 target_temp_reg_24_ ( .D(n2256), .CK(clk), .SN(rst_n), .Q(n6172), 
        .QN(target_temp[24]) );
  DFFSX1 target_temp_reg_23_ ( .D(n2255), .CK(clk), .SN(rst_n), .Q(n6167), 
        .QN(target_temp[23]) );
  DFFSX1 target_temp_reg_21_ ( .D(n2253), .CK(clk), .SN(rst_n), .Q(n6215), 
        .QN(target_temp[21]) );
  DFFSX1 target_temp_reg_20_ ( .D(n2252), .CK(clk), .SN(rst_n), .Q(n6166), 
        .QN(target_temp[20]) );
  DFFSX1 target_temp_reg_19_ ( .D(n2251), .CK(clk), .SN(rst_n), .Q(n6205), 
        .QN(target_temp[19]) );
  DFFSX1 target_temp_reg_18_ ( .D(n2250), .CK(clk), .SN(rst_n), .Q(n6186), 
        .QN(target_temp[18]) );
  DFFSX1 target_temp_reg_17_ ( .D(n2249), .CK(clk), .SN(rst_n), .Q(n6187), 
        .QN(target_temp[17]) );
  DFFSX1 target_temp_reg_16_ ( .D(n2248), .CK(clk), .SN(rst_n), .Q(n6207), 
        .QN(target_temp[16]) );
  DFFSX1 target_temp_reg_15_ ( .D(n2247), .CK(clk), .SN(rst_n), .Q(n6209), 
        .QN(target_temp[15]) );
  DFFSX1 target_temp_reg_14_ ( .D(n2246), .CK(clk), .SN(rst_n), .Q(n6211), 
        .QN(target_temp[14]) );
  DFFSX1 target_temp_reg_13_ ( .D(n2245), .CK(clk), .SN(rst_n), .Q(n6183), 
        .QN(target_temp[13]) );
  DFFSX1 target_temp_reg_12_ ( .D(n2244), .CK(clk), .SN(rst_n), .Q(n6184), 
        .QN(target_temp[12]) );
  DFFSX1 target_temp_reg_11_ ( .D(n2243), .CK(clk), .SN(rst_n), .Q(n6213), 
        .QN(target_temp[11]) );
  DFFSX1 target_temp_reg_10_ ( .D(n2242), .CK(clk), .SN(rst_n), .Q(n6193), 
        .QN(target_temp[10]) );
  DFFSX1 target_temp_reg_8_ ( .D(n2240), .CK(clk), .SN(rst_n), .Q(n6181), .QN(
        target_temp[8]) );
  DFFSX1 target_temp_reg_7_ ( .D(n2239), .CK(clk), .SN(rst_n), .Q(n6180), .QN(
        target_temp[7]) );
  DFFSX1 target_temp_reg_6_ ( .D(n2238), .CK(clk), .SN(rst_n), .Q(n6214), .QN(
        target_temp[6]) );
  DFFSX1 target_temp_reg_5_ ( .D(n2237), .CK(clk), .SN(rst_n), .Q(n6179), .QN(
        target_temp[5]) );
  DFFSX1 target_temp_reg_4_ ( .D(n2236), .CK(clk), .SN(rst_n), .Q(n6196), .QN(
        target_temp[4]) );
  DFFSX1 target_temp_reg_0_ ( .D(n2232), .CK(clk), .SN(rst_n), .Q(n6203), .QN(
        target_temp[0]) );
  DFFSX1 w2_reg_2__31_ ( .D(n2231), .CK(clk), .SN(rst_n), .QN(w2[95]) );
  DFFSX1 w1_reg_8__31_ ( .D(n2135), .CK(clk), .SN(rst_n), .QN(w1[287]) );
  DFFSX1 w1_reg_8__30_ ( .D(n2131), .CK(clk), .SN(rst_n), .QN(w1[286]) );
  DFFSX1 w1_reg_8__29_ ( .D(n2127), .CK(clk), .SN(rst_n), .QN(w1[285]) );
  DFFSX1 w1_reg_8__28_ ( .D(n2123), .CK(clk), .SN(rst_n), .QN(w1[284]) );
  DFFSX1 w1_reg_8__27_ ( .D(n2119), .CK(clk), .SN(rst_n), .QN(w1[283]) );
  DFFSX1 w1_reg_8__26_ ( .D(n2115), .CK(clk), .SN(rst_n), .QN(w1[282]) );
  DFFSX1 w1_reg_8__25_ ( .D(n2111), .CK(clk), .SN(rst_n), .QN(w1[281]) );
  DFFSX1 w1_reg_8__24_ ( .D(n2107), .CK(clk), .SN(rst_n), .QN(w1[280]) );
  DFFSX1 w1_reg_8__23_ ( .D(n2103), .CK(clk), .SN(rst_n), .QN(w1[279]) );
  DFFSX1 w1_reg_8__22_ ( .D(n2099), .CK(clk), .SN(rst_n), .QN(w1[278]) );
  DFFSX1 w1_reg_8__21_ ( .D(n2095), .CK(clk), .SN(rst_n), .QN(w1[277]) );
  DFFSX1 w1_reg_8__20_ ( .D(n2091), .CK(clk), .SN(rst_n), .QN(w1[276]) );
  DFFSX1 w1_reg_8__19_ ( .D(n2087), .CK(clk), .SN(rst_n), .QN(w1[275]) );
  DFFSX1 w1_reg_8__18_ ( .D(n2083), .CK(clk), .SN(rst_n), .QN(w1[274]) );
  DFFSX1 w1_reg_8__17_ ( .D(n2079), .CK(clk), .SN(rst_n), .QN(w1[273]) );
  DFFSX1 w1_reg_8__16_ ( .D(n2075), .CK(clk), .SN(rst_n), .QN(w1[272]) );
  DFFSX1 w1_reg_8__15_ ( .D(n2071), .CK(clk), .SN(rst_n), .QN(w1[271]) );
  DFFSX1 w1_reg_8__14_ ( .D(n2067), .CK(clk), .SN(rst_n), .QN(w1[270]) );
  DFFSX1 w1_reg_8__13_ ( .D(n2063), .CK(clk), .SN(rst_n), .QN(w1[269]) );
  DFFSX1 w1_reg_8__12_ ( .D(n2059), .CK(clk), .SN(rst_n), .QN(w1[268]) );
  DFFSX1 w1_reg_8__10_ ( .D(n2051), .CK(clk), .SN(rst_n), .QN(w1[266]) );
  DFFSX1 w1_reg_8__9_ ( .D(n2047), .CK(clk), .SN(rst_n), .QN(w1[265]) );
  DFFSX1 w1_reg_8__8_ ( .D(n2043), .CK(clk), .SN(rst_n), .QN(w1[264]) );
  DFFSX1 w1_reg_8__7_ ( .D(n2039), .CK(clk), .SN(rst_n), .QN(w1[263]) );
  DFFSX1 w1_reg_8__6_ ( .D(n2035), .CK(clk), .SN(rst_n), .QN(w1[262]) );
  DFFSX1 w1_reg_8__5_ ( .D(n2031), .CK(clk), .SN(rst_n), .QN(w1[261]) );
  DFFSX1 w1_reg_8__4_ ( .D(n2027), .CK(clk), .SN(rst_n), .QN(w1[260]) );
  DFFSX1 w1_reg_8__3_ ( .D(n2023), .CK(clk), .SN(rst_n), .QN(w1[259]) );
  DFFSX1 w1_reg_8__2_ ( .D(n2019), .CK(clk), .SN(rst_n), .QN(w1[258]) );
  DFFSX1 w1_reg_8__1_ ( .D(n2015), .CK(clk), .SN(rst_n), .QN(w1[257]) );
  DFFSX1 w1_reg_8__0_ ( .D(n2011), .CK(clk), .SN(rst_n), .QN(w1[256]) );
  DFFSX1 w1_reg_5__31_ ( .D(n2004), .CK(clk), .SN(rst_n), .QN(w1[191]) );
  DFFSX1 w1_reg_4__30_ ( .D(n2003), .CK(clk), .SN(rst_n), .QN(w1[158]) );
  DFFSX1 w1_reg_4__29_ ( .D(n1999), .CK(clk), .SN(rst_n), .QN(w1[157]) );
  DFFSX1 w1_reg_5__29_ ( .D(n1996), .CK(clk), .SN(rst_n), .QN(w1[189]) );
  DFFSX1 w1_reg_4__28_ ( .D(n1995), .CK(clk), .SN(rst_n), .QN(w1[156]) );
  DFFSX1 w1_reg_5__28_ ( .D(n1992), .CK(clk), .SN(rst_n), .QN(w1[188]) );
  DFFSX1 w1_reg_4__27_ ( .D(n1991), .CK(clk), .SN(rst_n), .QN(w1[155]) );
  DFFSX1 w1_reg_4__26_ ( .D(n1987), .CK(clk), .SN(rst_n), .QN(w1[154]) );
  DFFSX1 w1_reg_4__25_ ( .D(n1983), .CK(clk), .SN(rst_n), .QN(w1[153]) );
  DFFSX1 w1_reg_4__24_ ( .D(n1979), .CK(clk), .SN(rst_n), .QN(w1[152]) );
  DFFSX1 w1_reg_5__24_ ( .D(n1976), .CK(clk), .SN(rst_n), .QN(w1[184]) );
  DFFSX1 w1_reg_4__23_ ( .D(n1975), .CK(clk), .SN(rst_n), .QN(w1[151]) );
  DFFSX1 w1_reg_5__23_ ( .D(n1972), .CK(clk), .SN(rst_n), .QN(w1[183]) );
  DFFSX1 w1_reg_4__22_ ( .D(n1971), .CK(clk), .SN(rst_n), .QN(w1[150]) );
  DFFSX1 w1_reg_5__22_ ( .D(n1968), .CK(clk), .SN(rst_n), .QN(w1[182]) );
  DFFSX1 w1_reg_4__21_ ( .D(n1967), .CK(clk), .SN(rst_n), .QN(w1[149]) );
  DFFSX1 w1_reg_5__21_ ( .D(n1964), .CK(clk), .SN(rst_n), .QN(w1[181]) );
  DFFSX1 w1_reg_4__20_ ( .D(n1963), .CK(clk), .SN(rst_n), .QN(w1[148]) );
  DFFSX1 w1_reg_5__20_ ( .D(n1960), .CK(clk), .SN(rst_n), .QN(w1[180]) );
  DFFSX1 w1_reg_4__18_ ( .D(n1955), .CK(clk), .SN(rst_n), .QN(w1[146]) );
  DFFSX1 w1_reg_4__17_ ( .D(n1951), .CK(clk), .SN(rst_n), .QN(w1[145]) );
  DFFSX1 w1_reg_5__17_ ( .D(n1948), .CK(clk), .SN(rst_n), .QN(w1[177]) );
  DFFSX1 w1_reg_6__16_ ( .D(n1945), .CK(clk), .SN(rst_n), .QN(w1[208]) );
  DFFSX1 w1_reg_4__15_ ( .D(n1943), .CK(clk), .SN(rst_n), .QN(w1[143]) );
  DFFSX1 w1_reg_5__15_ ( .D(n1940), .CK(clk), .SN(rst_n), .QN(w1[175]) );
  DFFSX1 w1_reg_4__14_ ( .D(n1939), .CK(clk), .SN(rst_n), .QN(w1[142]) );
  DFFSX1 w1_reg_5__14_ ( .D(n1936), .CK(clk), .SN(rst_n), .QN(w1[174]) );
  DFFSX1 w1_reg_4__13_ ( .D(n1935), .CK(clk), .SN(rst_n), .QN(w1[141]) );
  DFFSX1 w1_reg_4__12_ ( .D(n1931), .CK(clk), .SN(rst_n), .QN(w1[140]) );
  DFFSX1 w1_reg_5__12_ ( .D(n1928), .CK(clk), .SN(rst_n), .QN(w1[172]) );
  DFFSX1 w1_reg_4__11_ ( .D(n1927), .CK(clk), .SN(rst_n), .QN(w1[139]) );
  DFFSX1 w1_reg_5__11_ ( .D(n1924), .CK(clk), .SN(rst_n), .QN(w1[171]) );
  DFFSX1 w1_reg_4__7_ ( .D(n1911), .CK(clk), .SN(rst_n), .QN(w1[135]) );
  DFFSX1 w1_reg_5__7_ ( .D(n1908), .CK(clk), .SN(rst_n), .QN(w1[167]) );
  DFFSX1 w1_reg_4__6_ ( .D(n1907), .CK(clk), .SN(rst_n), .QN(w1[134]) );
  DFFSX1 w1_reg_5__6_ ( .D(n1904), .CK(clk), .SN(rst_n), .QN(w1[166]) );
  DFFSX1 w1_reg_4__5_ ( .D(n1903), .CK(clk), .SN(rst_n), .QN(w1[133]) );
  DFFSX1 w1_reg_5__5_ ( .D(n1900), .CK(clk), .SN(rst_n), .QN(w1[165]) );
  DFFSX1 w1_reg_4__4_ ( .D(n1899), .CK(clk), .SN(rst_n), .QN(w1[132]) );
  DFFSX1 w1_reg_5__4_ ( .D(n1896), .CK(clk), .SN(rst_n), .QN(w1[164]) );
  DFFSX1 w1_reg_4__3_ ( .D(n1895), .CK(clk), .SN(rst_n), .QN(w1[131]) );
  DFFSX1 w1_reg_5__3_ ( .D(n1892), .CK(clk), .SN(rst_n), .QN(w1[163]) );
  DFFSX1 w1_reg_4__2_ ( .D(n1891), .CK(clk), .SN(rst_n), .QN(w1[130]) );
  DFFSX1 w1_reg_4__1_ ( .D(n1887), .CK(clk), .SN(rst_n), .QN(w1[129]) );
  DFFSX1 w1_reg_5__1_ ( .D(n1884), .CK(clk), .SN(rst_n), .QN(w1[161]) );
  DFFSX1 w1_reg_4__0_ ( .D(n1883), .CK(clk), .SN(rst_n), .QN(w1[128]) );
  DFFSX1 w1_reg_0__31_ ( .D(n1879), .CK(clk), .SN(rst_n), .QN(w1[31]) );
  DFFSX1 w1_reg_2__31_ ( .D(n1877), .CK(clk), .SN(rst_n), .QN(w1[95]) );
  DFFSX1 w1_reg_1__31_ ( .D(n1876), .CK(clk), .SN(rst_n), .QN(w1[63]) );
  DFFSX1 w1_reg_0__30_ ( .D(n1875), .CK(clk), .SN(rst_n), .QN(w1[30]) );
  DFFSX1 w1_reg_2__30_ ( .D(n1873), .CK(clk), .SN(rst_n), .QN(w1[94]) );
  DFFSX1 w1_reg_1__30_ ( .D(n1872), .CK(clk), .SN(rst_n), .QN(w1[62]) );
  DFFSX1 w1_reg_2__29_ ( .D(n1869), .CK(clk), .SN(rst_n), .QN(w1[93]) );
  DFFSX1 w1_reg_0__28_ ( .D(n1867), .CK(clk), .SN(rst_n), .QN(w1[28]) );
  DFFSX1 w1_reg_2__28_ ( .D(n1865), .CK(clk), .SN(rst_n), .QN(w1[92]) );
  DFFSX1 w1_reg_1__28_ ( .D(n1864), .CK(clk), .SN(rst_n), .QN(w1[60]) );
  DFFSX1 w1_reg_2__27_ ( .D(n1861), .CK(clk), .SN(rst_n), .QN(w1[91]) );
  DFFSX1 w1_reg_0__26_ ( .D(n1859), .CK(clk), .SN(rst_n), .QN(w1[26]) );
  DFFSX1 w1_reg_2__26_ ( .D(n1857), .CK(clk), .SN(rst_n), .QN(w1[90]) );
  DFFSX1 w1_reg_1__26_ ( .D(n1856), .CK(clk), .SN(rst_n), .QN(w1[58]) );
  DFFSX1 w1_reg_0__25_ ( .D(n1855), .CK(clk), .SN(rst_n), .QN(w1[25]) );
  DFFSX1 w1_reg_2__25_ ( .D(n1853), .CK(clk), .SN(rst_n), .QN(w1[89]) );
  DFFSX1 w1_reg_1__25_ ( .D(n1852), .CK(clk), .SN(rst_n), .QN(w1[57]) );
  DFFSX1 w1_reg_0__24_ ( .D(n1851), .CK(clk), .SN(rst_n), .QN(w1[24]) );
  DFFSX1 w1_reg_2__24_ ( .D(n1849), .CK(clk), .SN(rst_n), .QN(w1[88]) );
  DFFSX1 w1_reg_1__24_ ( .D(n1848), .CK(clk), .SN(rst_n), .QN(w1[56]) );
  DFFSX1 w1_reg_0__23_ ( .D(n1847), .CK(clk), .SN(rst_n), .QN(w1[23]) );
  DFFSX1 w1_reg_2__23_ ( .D(n1845), .CK(clk), .SN(rst_n), .QN(w1[87]) );
  DFFSX1 w1_reg_1__23_ ( .D(n1844), .CK(clk), .SN(rst_n), .QN(w1[55]) );
  DFFSX1 w1_reg_0__22_ ( .D(n1843), .CK(clk), .SN(rst_n), .QN(w1[22]) );
  DFFSX1 w1_reg_1__22_ ( .D(n1840), .CK(clk), .SN(rst_n), .QN(w1[54]) );
  DFFSX1 w1_reg_0__21_ ( .D(n1839), .CK(clk), .SN(rst_n), .QN(w1[21]) );
  DFFSX1 w1_reg_2__21_ ( .D(n1837), .CK(clk), .SN(rst_n), .QN(w1[85]) );
  DFFSX1 w1_reg_1__21_ ( .D(n1836), .CK(clk), .SN(rst_n), .QN(w1[53]) );
  DFFSX1 w1_reg_0__20_ ( .D(n1835), .CK(clk), .SN(rst_n), .QN(w1[20]) );
  DFFSX1 w1_reg_2__20_ ( .D(n1833), .CK(clk), .SN(rst_n), .QN(w1[84]) );
  DFFSX1 w1_reg_1__20_ ( .D(n1832), .CK(clk), .SN(rst_n), .QN(w1[52]) );
  DFFSX1 w1_reg_0__19_ ( .D(n1831), .CK(clk), .SN(rst_n), .QN(w1[19]) );
  DFFSX1 w1_reg_0__18_ ( .D(n1827), .CK(clk), .SN(rst_n), .QN(w1[18]) );
  DFFSX1 w1_reg_1__18_ ( .D(n1824), .CK(clk), .SN(rst_n), .QN(w1[50]) );
  DFFSX1 w1_reg_2__17_ ( .D(n1821), .CK(clk), .SN(rst_n), .QN(w1[81]) );
  DFFSX1 w1_reg_0__16_ ( .D(n1819), .CK(clk), .SN(rst_n), .QN(w1[16]) );
  DFFSX1 w1_reg_0__15_ ( .D(n1815), .CK(clk), .SN(rst_n), .QN(w1[15]) );
  DFFSX1 w1_reg_2__15_ ( .D(n1813), .CK(clk), .SN(rst_n), .QN(w1[79]) );
  DFFSX1 w1_reg_1__15_ ( .D(n1812), .CK(clk), .SN(rst_n), .QN(w1[47]) );
  DFFSX1 w1_reg_2__14_ ( .D(n1809), .CK(clk), .SN(rst_n), .QN(w1[78]) );
  DFFSX1 w1_reg_0__13_ ( .D(n1807), .CK(clk), .SN(rst_n), .QN(w1[13]) );
  DFFSX1 w1_reg_2__13_ ( .D(n1805), .CK(clk), .SN(rst_n), .QN(w1[77]) );
  DFFSX1 w1_reg_1__13_ ( .D(n1804), .CK(clk), .SN(rst_n), .QN(w1[45]) );
  DFFSX1 w1_reg_0__11_ ( .D(n1799), .CK(clk), .SN(rst_n), .QN(w1[11]) );
  DFFSX1 w1_reg_2__11_ ( .D(n1797), .CK(clk), .SN(rst_n), .QN(w1[75]) );
  DFFSX1 w1_reg_1__11_ ( .D(n1796), .CK(clk), .SN(rst_n), .QN(w1[43]) );
  DFFSX1 w1_reg_0__10_ ( .D(n1795), .CK(clk), .SN(rst_n), .QN(w1[10]) );
  DFFSX1 w1_reg_2__9_ ( .D(n1789), .CK(clk), .SN(rst_n), .QN(w1[73]) );
  DFFSX1 w1_reg_1__9_ ( .D(n1788), .CK(clk), .SN(rst_n), .QN(w1[41]) );
  DFFSX1 w1_reg_0__8_ ( .D(n1787), .CK(clk), .SN(rst_n), .QN(w1[8]) );
  DFFSX1 w1_reg_2__8_ ( .D(n1785), .CK(clk), .SN(rst_n), .QN(w1[72]) );
  DFFSX1 w1_reg_1__8_ ( .D(n1784), .CK(clk), .SN(rst_n), .QN(w1[40]) );
  DFFSX1 w1_reg_0__7_ ( .D(n1783), .CK(clk), .SN(rst_n), .QN(w1[7]) );
  DFFSX1 w1_reg_2__7_ ( .D(n1781), .CK(clk), .SN(rst_n), .QN(w1[71]) );
  DFFSX1 w1_reg_1__7_ ( .D(n1780), .CK(clk), .SN(rst_n), .QN(w1[39]) );
  DFFSX1 w1_reg_0__6_ ( .D(n1779), .CK(clk), .SN(rst_n), .QN(w1[6]) );
  DFFSX1 w1_reg_1__6_ ( .D(n1776), .CK(clk), .SN(rst_n), .QN(w1[38]) );
  DFFSX1 w1_reg_0__4_ ( .D(n1771), .CK(clk), .SN(rst_n), .QN(w1[4]) );
  DFFSX1 w1_reg_1__4_ ( .D(n1768), .CK(clk), .SN(rst_n), .QN(w1[36]) );
  DFFSX1 w1_reg_2__3_ ( .D(n1765), .CK(clk), .SN(rst_n), .QN(w1[67]) );
  DFFSX1 w1_reg_2__2_ ( .D(n1761), .CK(clk), .SN(rst_n), .QN(w1[66]) );
  DFFSX1 w1_reg_1__1_ ( .D(n1756), .CK(clk), .SN(rst_n), .QN(w1[33]) );
  DFFSX1 iter_reg_0_ ( .D(n1750), .CK(clk), .SN(rst_n), .QN(iter[0]) );
  DFFSX1 iter_reg_8_ ( .D(n1749), .CK(clk), .SN(rst_n), .QN(iter[8]) );
  DFFSX1 iter_reg_7_ ( .D(n1748), .CK(clk), .SN(rst_n), .Q(n26308) );
  DFFSX1 iter_reg_6_ ( .D(n1747), .CK(clk), .SN(rst_n), .QN(iter[6]) );
  DFFSX1 iter_reg_4_ ( .D(n1745), .CK(clk), .SN(rst_n), .QN(iter[4]) );
  DFFSX1 iter_reg_3_ ( .D(n1744), .CK(clk), .SN(rst_n), .Q(n26309) );
  DFFSX1 iter_reg_2_ ( .D(n1743), .CK(clk), .SN(rst_n), .QN(iter[2]) );
  DFFSX1 data_reg_3__31_ ( .D(n1741), .CK(clk), .SN(rst_n), .QN(data[127]) );
  DFFSX1 data_reg_3__30_ ( .D(n1740), .CK(clk), .SN(rst_n), .QN(data[126]) );
  DFFSX1 data_reg_3__29_ ( .D(n1739), .CK(clk), .SN(rst_n), .QN(data[125]) );
  DFFSX1 data_reg_3__28_ ( .D(n1738), .CK(clk), .SN(rst_n), .QN(data[124]) );
  DFFSX1 data_reg_3__27_ ( .D(n1737), .CK(clk), .SN(rst_n), .QN(data[123]) );
  DFFSX1 data_reg_3__26_ ( .D(n1736), .CK(clk), .SN(rst_n), .QN(data[122]) );
  DFFSX1 data_reg_3__25_ ( .D(n1735), .CK(clk), .SN(rst_n), .QN(data[121]) );
  DFFSX1 data_reg_3__24_ ( .D(n1734), .CK(clk), .SN(rst_n), .QN(data[120]) );
  DFFSX1 data_reg_3__23_ ( .D(n1733), .CK(clk), .SN(rst_n), .QN(data[119]) );
  DFFSX1 data_reg_2__31_ ( .D(n1709), .CK(clk), .SN(rst_n), .QN(data[95]) );
  DFFSX1 data_reg_2__30_ ( .D(n1708), .CK(clk), .SN(rst_n), .QN(data[94]) );
  DFFSX1 data_reg_2__29_ ( .D(n1707), .CK(clk), .SN(rst_n), .QN(data[93]) );
  DFFSX1 data_reg_2__28_ ( .D(n1706), .CK(clk), .SN(rst_n), .QN(data[92]) );
  DFFSX1 data_reg_2__27_ ( .D(n1705), .CK(clk), .SN(rst_n), .QN(data[91]) );
  DFFSX1 data_reg_2__26_ ( .D(n1704), .CK(clk), .SN(rst_n), .QN(data[90]) );
  DFFSX1 data_reg_2__25_ ( .D(n1703), .CK(clk), .SN(rst_n), .QN(data[89]) );
  DFFSX1 data_reg_2__24_ ( .D(n1702), .CK(clk), .SN(rst_n), .QN(data[88]) );
  DFFSX1 data_reg_2__23_ ( .D(n1701), .CK(clk), .SN(rst_n), .Q(n2986), .QN(
        data[87]) );
  DFFSX1 data_reg_1__31_ ( .D(n1677), .CK(clk), .SN(rst_n), .QN(data[63]) );
  DFFSX1 data_reg_1__30_ ( .D(n1676), .CK(clk), .SN(rst_n), .QN(data[62]) );
  DFFSX1 data_reg_1__29_ ( .D(n1675), .CK(clk), .SN(rst_n), .QN(data[61]) );
  DFFSX1 data_reg_1__28_ ( .D(n1674), .CK(clk), .SN(rst_n), .QN(data[60]) );
  DFFSX1 data_reg_1__27_ ( .D(n1673), .CK(clk), .SN(rst_n), .QN(data[59]) );
  DFFSX1 data_reg_1__26_ ( .D(n1672), .CK(clk), .SN(rst_n), .QN(data[58]) );
  DFFSX1 data_reg_1__25_ ( .D(n1671), .CK(clk), .SN(rst_n), .QN(data[57]) );
  DFFSX1 data_reg_1__24_ ( .D(n1670), .CK(clk), .SN(rst_n), .QN(data[56]) );
  DFFSX1 data_reg_1__23_ ( .D(n1669), .CK(clk), .SN(rst_n), .QN(data[55]) );
  DFFSX1 data_reg_0__31_ ( .D(n1645), .CK(clk), .SN(rst_n), .QN(data[31]) );
  DFFSX1 data_reg_0__30_ ( .D(n1644), .CK(clk), .SN(rst_n), .QN(data[30]) );
  DFFSX1 data_reg_0__29_ ( .D(n1643), .CK(clk), .SN(rst_n), .QN(data[29]) );
  DFFSX1 data_reg_0__28_ ( .D(n1642), .CK(clk), .SN(rst_n), .QN(data[28]) );
  DFFSX1 data_reg_0__27_ ( .D(n1641), .CK(clk), .SN(rst_n), .QN(data[27]) );
  DFFSX1 data_reg_0__26_ ( .D(n1640), .CK(clk), .SN(rst_n), .QN(data[26]) );
  DFFSX1 data_reg_0__25_ ( .D(n1639), .CK(clk), .SN(rst_n), .QN(data[25]) );
  DFFSX1 data_reg_0__24_ ( .D(n1638), .CK(clk), .SN(rst_n), .QN(data[24]) );
  DFFSX1 data_reg_0__23_ ( .D(n1637), .CK(clk), .SN(rst_n), .QN(data[23]) );
  DFFSX1 data_reg_0__22_ ( .D(n1636), .CK(clk), .SN(rst_n), .QN(data[22]) );
  DFFSX1 data_reg_0__21_ ( .D(n1635), .CK(clk), .SN(rst_n), .QN(data[21]) );
  DFFSX1 data_reg_0__20_ ( .D(n1634), .CK(clk), .SN(rst_n), .QN(data[20]) );
  DFFSX1 data_reg_0__19_ ( .D(n1633), .CK(clk), .SN(rst_n), .QN(data[19]) );
  DFFSX1 data_reg_0__18_ ( .D(n1632), .CK(clk), .SN(rst_n), .QN(data[18]) );
  DFFSX1 data_reg_0__17_ ( .D(n1631), .CK(clk), .SN(rst_n), .QN(data[17]) );
  DFFSX1 data_reg_0__16_ ( .D(n1630), .CK(clk), .SN(rst_n), .QN(data[16]) );
  DFFSX1 data_reg_0__15_ ( .D(n1629), .CK(clk), .SN(rst_n), .QN(data[15]) );
  DFFSX1 data_reg_0__14_ ( .D(n1628), .CK(clk), .SN(rst_n), .QN(data[14]) );
  DFFSX1 data_reg_0__13_ ( .D(n1627), .CK(clk), .SN(rst_n), .QN(data[13]) );
  DFFSX1 data_reg_0__12_ ( .D(n1626), .CK(clk), .SN(rst_n), .QN(data[12]) );
  DFFSX1 data_reg_0__11_ ( .D(n1625), .CK(clk), .SN(rst_n), .QN(data[11]) );
  DFFSX1 data_reg_0__10_ ( .D(n1624), .CK(clk), .SN(rst_n), .QN(data[10]) );
  DFFSX1 data_reg_0__9_ ( .D(n1623), .CK(clk), .SN(rst_n), .QN(data[9]) );
  DFFSX1 data_reg_0__8_ ( .D(n1622), .CK(clk), .SN(rst_n), .QN(data[8]) );
  DFFSX1 data_reg_0__7_ ( .D(n1621), .CK(clk), .SN(rst_n), .QN(data[7]) );
  DFFSX1 data_reg_0__6_ ( .D(n1620), .CK(clk), .SN(rst_n), .QN(data[6]) );
  DFFSX1 data_reg_0__5_ ( .D(n1619), .CK(clk), .SN(rst_n), .QN(data[5]) );
  DFFSX1 data_reg_0__4_ ( .D(n1618), .CK(clk), .SN(rst_n), .QN(data[4]) );
  DFFSX1 data_reg_0__3_ ( .D(n1617), .CK(clk), .SN(rst_n), .QN(data[3]) );
  DFFSX1 data_reg_0__2_ ( .D(n1616), .CK(clk), .SN(rst_n), .QN(data[2]) );
  DFFSX1 data_reg_0__1_ ( .D(n1615), .CK(clk), .SN(rst_n), .QN(data[1]) );
  DFFSX1 data_reg_0__0_ ( .D(n1614), .CK(clk), .SN(rst_n), .QN(data[0]) );
  CMPR42X1 M6_mult_x_15_U570 ( .A(M6_mult_x_15_n724), .B(M6_mult_x_15_n1159), 
        .C(M6_mult_x_15_n727), .D(M6_mult_x_15_n1183), .ICI(M6_mult_x_15_n1207), .S(M6_mult_x_15_n722), .ICO(M6_mult_x_15_n720), .CO(M6_mult_x_15_n721) );
  CMPR42X1 M6_mult_x_15_U568 ( .A(M6_mult_x_15_n719), .B(M6_mult_x_15_n1158), 
        .C(M6_mult_x_15_n720), .D(M6_mult_x_15_n1182), .ICI(M6_mult_x_15_n1206), .S(M6_mult_x_15_n717), .ICO(M6_mult_x_15_n715), .CO(M6_mult_x_15_n716) );
  CMPR42X1 M6_mult_x_15_U566 ( .A(M6_mult_x_15_n714), .B(M6_mult_x_15_n1157), 
        .C(M6_mult_x_15_n715), .D(M6_mult_x_15_n1181), .ICI(M6_mult_x_15_n1205), .S(M6_mult_x_15_n712), .ICO(M6_mult_x_15_n710), .CO(M6_mult_x_15_n711) );
  CMPR42X1 M6_mult_x_15_U560 ( .A(M6_mult_x_15_n1155), .B(M6_mult_x_15_n1203), 
        .C(M6_mult_x_15_n1179), .D(M6_mult_x_15_n700), .ICI(M6_mult_x_15_n703), 
        .S(M6_mult_x_15_n698), .ICO(M6_mult_x_15_n696), .CO(M6_mult_x_15_n697)
         );
  CMPR42X1 M6_mult_x_15_U557 ( .A(M6_mult_x_15_n1154), .B(M6_mult_x_15_n1178), 
        .C(M6_mult_x_15_n1202), .D(M6_mult_x_15_n693), .ICI(M6_mult_x_15_n696), 
        .S(M6_mult_x_15_n691), .ICO(M6_mult_x_15_n689), .CO(M6_mult_x_15_n690)
         );
  CMPR42X1 M6_mult_x_15_U555 ( .A(M6_mult_x_15_n688), .B(M6_mult_x_15_n1105), 
        .C(M6_mult_x_15_n694), .D(M6_mult_x_15_n1129), .ICI(M6_mult_x_15_n1153), .S(M6_mult_x_15_n686), .ICO(M6_mult_x_15_n684), .CO(M6_mult_x_15_n685) );
  CMPR42X1 M6_mult_x_15_U554 ( .A(M6_mult_x_15_n1201), .B(M6_mult_x_15_n1177), 
        .C(M6_mult_x_15_n692), .D(M6_mult_x_15_n689), .ICI(M6_mult_x_15_n686), 
        .S(M6_mult_x_15_n683), .ICO(M6_mult_x_15_n681), .CO(M6_mult_x_15_n682)
         );
  CMPR42X1 M6_mult_x_15_U552 ( .A(M6_mult_x_15_n680), .B(M6_mult_x_15_n1104), 
        .C(M6_mult_x_15_n684), .D(M6_mult_x_15_n1128), .ICI(M6_mult_x_15_n1176), .S(M6_mult_x_15_n678), .ICO(M6_mult_x_15_n676), .CO(M6_mult_x_15_n677) );
  CMPR42X1 M6_mult_x_15_U551 ( .A(M6_mult_x_15_n1152), .B(M6_mult_x_15_n1200), 
        .C(M6_mult_x_15_n685), .D(M6_mult_x_15_n681), .ICI(M6_mult_x_15_n678), 
        .S(M6_mult_x_15_n675), .ICO(M6_mult_x_15_n673), .CO(M6_mult_x_15_n674)
         );
  CMPR42X1 M6_mult_x_15_U549 ( .A(M6_mult_x_15_n672), .B(M6_mult_x_15_n1103), 
        .C(M6_mult_x_15_n676), .D(M6_mult_x_15_n1127), .ICI(M6_mult_x_15_n1199), .S(M6_mult_x_15_n670), .ICO(M6_mult_x_15_n668), .CO(M6_mult_x_15_n669) );
  CMPR42X1 M6_mult_x_15_U548 ( .A(M6_mult_x_15_n1151), .B(M6_mult_x_15_n1175), 
        .C(M6_mult_x_15_n677), .D(M6_mult_x_15_n673), .ICI(M6_mult_x_15_n670), 
        .S(M6_mult_x_15_n667), .ICO(M6_mult_x_15_n665), .CO(M6_mult_x_15_n666)
         );
  CMPR42X1 M6_mult_x_15_U544 ( .A(M6_mult_x_15_n1150), .B(M6_mult_x_15_n1198), 
        .C(M6_mult_x_15_n669), .D(M6_mult_x_15_n665), .ICI(M6_mult_x_15_n660), 
        .S(M6_mult_x_15_n657), .ICO(M6_mult_x_15_n655), .CO(M6_mult_x_15_n656)
         );
  CMPR42X1 M6_mult_x_15_U541 ( .A(M6_mult_x_15_n1101), .B(M6_mult_x_15_n1149), 
        .C(M6_mult_x_15_n1125), .D(M6_mult_x_15_n658), .ICI(M6_mult_x_15_n1197), .S(M6_mult_x_15_n650), .ICO(M6_mult_x_15_n648), .CO(M6_mult_x_15_n649) );
  CMPR42X1 M6_mult_x_15_U536 ( .A(M6_mult_x_15_n1124), .B(M6_mult_x_15_n642), 
        .C(M6_mult_x_15_n649), .D(M6_mult_x_15_n645), .ICI(M6_mult_x_15_n640), 
        .S(M6_mult_x_15_n637), .ICO(M6_mult_x_15_n635), .CO(M6_mult_x_15_n636)
         );
  CMPR42X1 M6_mult_x_15_U534 ( .A(M6_mult_x_15_n634), .B(M6_mult_x_15_n1051), 
        .C(M6_mult_x_15_n643), .D(M6_mult_x_15_n1075), .ICI(M6_mult_x_15_n1099), .S(M6_mult_x_15_n632), .ICO(M6_mult_x_15_n630), .CO(M6_mult_x_15_n631) );
  CMPR42X1 M6_mult_x_15_U533 ( .A(M6_mult_x_15_n1147), .B(M6_mult_x_15_n1123), 
        .C(M6_mult_x_15_n1171), .D(M6_mult_x_15_n641), .ICI(M6_mult_x_15_n632), 
        .S(M6_mult_x_15_n629), .ICO(M6_mult_x_15_n627), .CO(M6_mult_x_15_n628)
         );
  CMPR42X1 M6_mult_x_15_U532 ( .A(M6_mult_x_15_n1195), .B(M6_mult_x_15_n638), 
        .C(M6_mult_x_15_n639), .D(M6_mult_x_15_n629), .ICI(M6_mult_x_15_n635), 
        .S(M6_mult_x_15_n626), .ICO(M6_mult_x_15_n624), .CO(M6_mult_x_15_n625)
         );
  CMPR42X1 M6_mult_x_15_U530 ( .A(M6_mult_x_15_n623), .B(M6_mult_x_15_n1050), 
        .C(M6_mult_x_15_n630), .D(M6_mult_x_15_n1074), .ICI(M6_mult_x_15_n1098), .S(M6_mult_x_15_n621), .ICO(M6_mult_x_15_n619), .CO(M6_mult_x_15_n620) );
  CMPR42X1 M6_mult_x_15_U526 ( .A(M6_mult_x_15_n612), .B(M6_mult_x_15_n1049), 
        .C(M6_mult_x_15_n619), .D(M6_mult_x_15_n1073), .ICI(M6_mult_x_15_n1097), .S(M6_mult_x_15_n610), .ICO(M6_mult_x_15_n608), .CO(M6_mult_x_15_n609) );
  CMPR42X1 M6_mult_x_15_U524 ( .A(M6_mult_x_15_n620), .B(M6_mult_x_15_n610), 
        .C(M6_mult_x_15_n617), .D(M6_mult_x_15_n607), .ICI(M6_mult_x_15_n613), 
        .S(M6_mult_x_15_n604), .ICO(M6_mult_x_15_n602), .CO(M6_mult_x_15_n603)
         );
  CMPR42X1 M6_mult_x_15_U522 ( .A(M6_mult_x_15_n601), .B(M6_mult_x_15_n1048), 
        .C(M6_mult_x_15_n1072), .D(M6_mult_x_15_n1120), .ICI(M6_mult_x_15_n608), .S(M6_mult_x_15_n599), .ICO(M6_mult_x_15_n597), .CO(M6_mult_x_15_n598) );
  CMPR42X1 M6_mult_x_15_U521 ( .A(M6_mult_x_15_n1192), .B(M6_mult_x_15_n1096), 
        .C(M6_mult_x_15_n1144), .D(M6_mult_x_15_n1168), .ICI(M6_mult_x_15_n609), .S(M6_mult_x_15_n596), .ICO(M6_mult_x_15_n594), .CO(M6_mult_x_15_n595) );
  CMPR42X1 M6_mult_x_15_U520 ( .A(M6_mult_x_15_n605), .B(M6_mult_x_15_n599), 
        .C(M6_mult_x_15_n606), .D(M6_mult_x_15_n596), .ICI(M6_mult_x_15_n602), 
        .S(M6_mult_x_15_n593), .ICO(M6_mult_x_15_n591), .CO(M6_mult_x_15_n592)
         );
  CMPR42X1 M6_mult_x_15_U518 ( .A(M6_mult_x_15_n1047), .B(M6_mult_x_15_n590), 
        .C(M6_mult_x_15_n1095), .D(M6_mult_x_15_n1191), .ICI(M6_mult_x_15_n594), .S(M6_mult_x_15_n588), .ICO(M6_mult_x_15_n586), .CO(M6_mult_x_15_n587) );
  CMPR42X1 M6_mult_x_15_U517 ( .A(M6_mult_x_15_n1071), .B(M6_mult_x_15_n597), 
        .C(M6_mult_x_15_n1119), .D(M6_mult_x_15_n1143), .ICI(M6_mult_x_15_n598), .S(M6_mult_x_15_n585), .ICO(M6_mult_x_15_n583), .CO(M6_mult_x_15_n584) );
  CMPR42X1 M6_mult_x_15_U514 ( .A(M6_mult_x_15_n589), .B(M6_mult_x_15_n579), 
        .C(M6_mult_x_15_n1046), .D(M6_mult_x_15_n1118), .ICI(M6_mult_x_15_n583), .S(M6_mult_x_15_n577), .ICO(M6_mult_x_15_n575), .CO(M6_mult_x_15_n576) );
  CMPR42X1 M6_mult_x_15_U510 ( .A(M6_mult_x_15_n578), .B(M6_mult_x_15_n1045), 
        .C(M6_mult_x_15_n568), .D(M6_mult_x_15_n1093), .ICI(M6_mult_x_15_n575), 
        .S(M6_mult_x_15_n566), .ICO(M6_mult_x_15_n564), .CO(M6_mult_x_15_n565)
         );
  CMPR42X1 M6_mult_x_15_U508 ( .A(M6_mult_x_15_n576), .B(M6_mult_x_15_n566), 
        .C(M6_mult_x_15_n573), .D(M6_mult_x_15_n563), .ICI(M6_mult_x_15_n569), 
        .S(M6_mult_x_15_n560), .ICO(M6_mult_x_15_n558), .CO(M6_mult_x_15_n559)
         );
  CMPR42X1 M6_mult_x_15_U505 ( .A(M6_mult_x_15_n1068), .B(M6_mult_x_15_n1092), 
        .C(M6_mult_x_15_n564), .D(M6_mult_x_15_n1116), .ICI(M6_mult_x_15_n565), 
        .S(M6_mult_x_15_n552), .ICO(M6_mult_x_15_n550), .CO(M6_mult_x_15_n551)
         );
  CMPR42X1 M6_mult_x_15_U502 ( .A(M6_mult_x_15_n546), .B(M6_mult_x_15_n1020), 
        .C(M6_mult_x_15_n556), .D(M6_mult_x_15_n1043), .ICI(M6_mult_x_15_n1091), .S(M6_mult_x_15_n544), .ICO(M6_mult_x_15_n542), .CO(M6_mult_x_15_n543) );
  CMPR42X1 M6_mult_x_15_U498 ( .A(n26495), .B(M6_mult_x_15_n545), .C(
        M6_mult_x_15_n1019), .D(M6_mult_x_15_n1066), .ICI(M6_mult_x_15_n1138), 
        .S(M6_mult_x_15_n534), .ICO(M6_mult_x_15_n532), .CO(M6_mult_x_15_n533)
         );
  CMPR42X1 M6_mult_x_15_U497 ( .A(M6_mult_x_15_n542), .B(M6_mult_x_15_n1042), 
        .C(M6_mult_x_15_n1090), .D(M6_mult_x_15_n1114), .ICI(M6_mult_x_15_n543), .S(M6_mult_x_15_n531), .ICO(M6_mult_x_15_n529), .CO(M6_mult_x_15_n530) );
  CMPR42X1 M6_mult_x_15_U496 ( .A(M6_mult_x_15_n539), .B(M6_mult_x_15_n534), 
        .C(M6_mult_x_15_n531), .D(M6_mult_x_15_n540), .ICI(M6_mult_x_15_n536), 
        .S(M6_mult_x_15_n528), .ICO(M6_mult_x_15_n526), .CO(M6_mult_x_15_n527)
         );
  CMPR42X1 M6_mult_x_15_U492 ( .A(M6_mult_x_15_n529), .B(M6_mult_x_15_n533), 
        .C(M6_mult_x_15_n530), .D(M6_mult_x_15_n521), .ICI(M6_mult_x_15_n526), 
        .S(M6_mult_x_15_n518), .ICO(M6_mult_x_15_n516), .CO(M6_mult_x_15_n517)
         );
  CMPR42X1 M6_mult_x_15_U489 ( .A(M6_mult_x_15_n519), .B(M6_mult_x_15_n515), 
        .C(M6_mult_x_15_n520), .D(M6_mult_x_15_n512), .ICI(M6_mult_x_15_n516), 
        .S(M6_mult_x_15_n509), .ICO(M6_mult_x_15_n507), .CO(M6_mult_x_15_n508)
         );
  CMPR42X1 M6_mult_x_15_U486 ( .A(M6_mult_x_15_n1016), .B(M6_mult_x_15_n1111), 
        .C(M6_mult_x_15_n1063), .D(M6_mult_x_15_n1087), .ICI(M6_mult_x_15_n510), .S(M6_mult_x_15_n503), .ICO(M6_mult_x_15_n501), .CO(M6_mult_x_15_n502) );
  CMPR42X1 M6_mult_x_15_U485 ( .A(M6_mult_x_15_n505), .B(M6_mult_x_15_n514), 
        .C(M6_mult_x_15_n503), .D(M6_mult_x_15_n511), .ICI(M6_mult_x_15_n507), 
        .S(M6_mult_x_15_n500), .ICO(M6_mult_x_15_n498), .CO(M6_mult_x_15_n499)
         );
  CMPR42X1 M6_mult_x_15_U482 ( .A(M6_mult_x_15_n1110), .B(M6_mult_x_15_n1038), 
        .C(M6_mult_x_15_n504), .D(M6_mult_x_15_n1086), .ICI(M6_mult_x_15_n501), 
        .S(M6_mult_x_15_n494), .ICO(M6_mult_x_15_n492), .CO(M6_mult_x_15_n493)
         );
  CMPR42X1 M6_mult_x_15_U479 ( .A(M6_mult_x_15_n488), .B(M6_mult_x_15_n1014), 
        .C(M6_mult_x_15_n1037), .D(M6_mult_x_15_n495), .ICI(M6_mult_x_15_n1085), .S(M6_mult_x_15_n486), .ICO(M6_mult_x_15_n484), .CO(M6_mult_x_15_n485) );
  CMPR42X1 M6_mult_x_15_U476 ( .A(n26492), .B(M6_mult_x_15_n487), .C(
        M6_mult_x_15_n1013), .D(M6_mult_x_15_n1084), .ICI(M6_mult_x_15_n1036), 
        .S(M6_mult_x_15_n479), .ICO(M6_mult_x_15_n477), .CO(M6_mult_x_15_n478)
         );
  CMPR42X1 M6_mult_x_15_U470 ( .A(M6_mult_x_15_n470), .B(M6_mult_x_15_n1034), 
        .C(M6_mult_x_15_n466), .D(M6_mult_x_15_n471), .ICI(M6_mult_x_15_n467), 
        .S(M6_mult_x_15_n463), .ICO(M6_mult_x_15_n461), .CO(M6_mult_x_15_n462)
         );
  CMPR42X1 M6_mult_x_15_U467 ( .A(M6_mult_x_15_n1010), .B(M6_mult_x_15_n1033), 
        .C(M6_mult_x_15_n459), .D(M6_mult_x_15_n465), .ICI(M6_mult_x_15_n461), 
        .S(M6_mult_x_15_n457), .ICO(M6_mult_x_15_n455), .CO(M6_mult_x_15_n456)
         );
  CMPR42X1 M6_mult_x_15_U464 ( .A(M6_mult_x_15_n1056), .B(M6_mult_x_15_n458), 
        .C(M6_mult_x_15_n453), .D(M6_mult_x_15_n1032), .ICI(M6_mult_x_15_n455), 
        .S(M6_mult_x_15_n451), .ICO(M6_mult_x_15_n449), .CO(M6_mult_x_15_n450)
         );
  CMPR42X1 M6_mult_x_15_U462 ( .A(M6_mult_x_15_n448), .B(M6_mult_x_15_n1031), 
        .C(M6_mult_x_15_n1008), .D(M6_mult_x_15_n452), .ICI(M6_mult_x_15_n449), 
        .S(M6_mult_x_15_n446), .ICO(M6_mult_x_15_n444), .CO(M6_mult_x_15_n445)
         );
  CMPR42X1 M6_mult_x_15_U460 ( .A(n26490), .B(M6_mult_x_15_n447), .C(
        M6_mult_x_15_n1030), .D(M6_mult_x_15_n1007), .ICI(M6_mult_x_15_n444), 
        .S(M6_mult_x_15_n442), .ICO(M6_mult_x_15_n440), .CO(M6_mult_x_15_n441)
         );
  CMPR42X1 M6_mult_x_15_U458 ( .A(n11074), .B(n26490), .C(M6_mult_x_15_n1029), 
        .D(M6_mult_x_15_n1006), .ICI(M6_mult_x_15_n440), .S(M6_mult_x_15_n438), 
        .ICO(M6_mult_x_15_n436), .CO(M6_mult_x_15_n437) );
  OAI21XL M2_U3_U1_UEN1_2_4_0 ( .A0(n25984), .A1(n26204), .B0(
        M2_U3_U1_enc_tree_2__3__24_), .Y(M2_U3_U1_enc_tree_2__4__16_) );
  OAI21XL M2_U3_U1_UEN1_1_4_0 ( .A0(M2_U3_U1_enc_tree_1__3__8_), .A1(n26205), 
        .B0(M2_U3_U1_enc_tree_1__3__24_), .Y(M2_U3_U1_enc_tree_1__4__16_) );
  OAI21XL M2_U3_U1_UEN1_1_2_3 ( .A0(M2_U3_U1_enc_tree_1__1__26_), .A1(
        M2_U3_U1_or2_inv_1__28_), .B0(M2_U3_U1_enc_tree_1__1__30_), .Y(
        M2_U3_U1_enc_tree_1__2__28_) );
  OAI21XL M2_U3_U1_UEN1_1_2_2 ( .A0(M2_U3_U1_enc_tree_1__1__18_), .A1(
        M2_U3_U1_or2_inv_1__20_), .B0(M2_U3_U1_enc_tree_1__1__22_), .Y(
        M2_U3_U1_enc_tree_1__2__20_) );
  OAI21XL M2_U3_U1_UEN1_1_2_1 ( .A0(M2_U3_U1_enc_tree_1__1__10_), .A1(
        M2_U3_U1_or2_inv_1__12_), .B0(M2_U3_U1_enc_tree_1__1__14_), .Y(
        M2_U3_U1_enc_tree_1__2__12_) );
  OAI21XL M2_U3_U1_UEN1_0_4_0 ( .A0(M2_U3_U1_enc_tree_0__3__8_), .A1(n26207), 
        .B0(M2_U3_U1_enc_tree_0__3__24_), .Y(M2_U3_U1_enc_tree_0__4__16_) );
  OAI21XL M2_U3_U1_UEN1_0_2_3 ( .A0(M2_U3_U1_enc_tree_0__1__26_), .A1(
        M2_U3_U1_or2_inv_0__28_), .B0(M2_U3_U1_enc_tree_0__1__30_), .Y(
        M2_U3_U1_enc_tree_0__2__28_) );
  OAI21XL M2_U3_U1_UEN1_0_2_2 ( .A0(M2_U3_U1_enc_tree_0__1__18_), .A1(
        M2_U3_U1_or2_inv_0__20_), .B0(M2_U3_U1_enc_tree_0__1__22_), .Y(
        M2_U3_U1_enc_tree_0__2__20_) );
  OAI21XL M2_U3_U1_UEN1_0_2_1 ( .A0(M2_U3_U1_enc_tree_0__1__10_), .A1(
        M2_U3_U1_or2_tree_0__1__12_), .B0(M2_U3_U1_enc_tree_0__1__14_), .Y(
        M2_U3_U1_enc_tree_0__2__12_) );
  OAI21XL M1_U3_U1_UEN1_2_4_0 ( .A0(n25987), .A1(n26199), .B0(
        M1_U3_U1_enc_tree_2__3__24_), .Y(M1_U3_U1_enc_tree_2__4__16_) );
  OAI21XL M1_U3_U1_UEN1_1_4_0 ( .A0(M1_U3_U1_enc_tree_1__3__8_), .A1(n26210), 
        .B0(M1_U3_U1_enc_tree_1__3__24_), .Y(M1_U3_U1_enc_tree_1__4__16_) );
  OAI21XL M1_U3_U1_UEN1_1_2_3 ( .A0(M1_U3_U1_enc_tree_1__1__26_), .A1(
        M1_U3_U1_or2_inv_1__28_), .B0(M1_U3_U1_enc_tree_1__1__30_), .Y(
        M1_U3_U1_enc_tree_1__2__28_) );
  OAI21XL M1_U3_U1_UEN1_1_2_2 ( .A0(M1_U3_U1_enc_tree_1__1__18_), .A1(
        M1_U3_U1_or2_inv_1__20_), .B0(M1_U3_U1_enc_tree_1__1__22_), .Y(
        M1_U3_U1_enc_tree_1__2__20_) );
  OAI21XL M1_U3_U1_UEN1_1_2_1 ( .A0(M1_U3_U1_enc_tree_1__1__10_), .A1(
        M1_U3_U1_or2_inv_1__12_), .B0(M1_U3_U1_enc_tree_1__1__14_), .Y(
        M1_U3_U1_enc_tree_1__2__12_) );
  OAI21XL M1_U3_U1_UEN1_0_4_0 ( .A0(M1_U3_U1_enc_tree_0__3__8_), .A1(n26209), 
        .B0(M1_U3_U1_enc_tree_0__3__24_), .Y(M1_U3_U1_enc_tree_0__4__16_) );
  OAI21XL M1_U3_U1_UEN1_0_2_3 ( .A0(M1_U3_U1_enc_tree_0__1__26_), .A1(
        M1_U3_U1_or2_inv_0__28_), .B0(M1_U3_U1_enc_tree_0__1__30_), .Y(
        M1_U3_U1_enc_tree_0__2__28_) );
  OAI21XL M1_U3_U1_UEN1_0_2_2 ( .A0(M1_U3_U1_enc_tree_0__1__18_), .A1(
        M1_U3_U1_or2_inv_0__20_), .B0(M1_U3_U1_enc_tree_0__1__22_), .Y(
        M1_U3_U1_enc_tree_0__2__20_) );
  OAI21XL M1_U3_U1_UEN1_0_2_1 ( .A0(M1_U3_U1_enc_tree_0__1__10_), .A1(
        M1_U3_U1_or2_tree_0__1__12_), .B0(M1_U3_U1_enc_tree_0__1__14_), .Y(
        M1_U3_U1_enc_tree_0__2__12_) );
  OAI21XL M2_U4_U1_UEN1_2_4_0 ( .A0(n25989), .A1(n26197), .B0(
        M2_U4_U1_enc_tree_2__3__24_), .Y(M2_U4_U1_enc_tree_2__4__16_) );
  OAI21XL M2_U4_U1_UEN1_1_4_0 ( .A0(M2_U4_U1_enc_tree_1__3__8_), .A1(n26153), 
        .B0(M2_U4_U1_enc_tree_1__3__24_), .Y(M2_U4_U1_enc_tree_1__4__16_) );
  OAI21XL M2_U4_U1_UEN1_1_2_3 ( .A0(M2_U4_U1_enc_tree_1__1__26_), .A1(
        M2_U4_U1_or2_inv_1__28_), .B0(M2_U4_U1_enc_tree_1__1__30_), .Y(
        M2_U4_U1_enc_tree_1__2__28_) );
  OAI21XL M2_U4_U1_UEN1_1_2_2 ( .A0(M2_U4_U1_enc_tree_1__1__18_), .A1(
        M2_U4_U1_or2_inv_1__20_), .B0(M2_U4_U1_enc_tree_1__1__22_), .Y(
        M2_U4_U1_enc_tree_1__2__20_) );
  OAI21XL M2_U4_U1_UEN1_1_2_1 ( .A0(M2_U4_U1_enc_tree_1__1__10_), .A1(
        M2_U4_U1_or2_inv_1__12_), .B0(M2_U4_U1_enc_tree_1__1__14_), .Y(
        M2_U4_U1_enc_tree_1__2__12_) );
  OAI21XL M2_U4_U1_UEN1_0_4_0 ( .A0(M2_U4_U1_enc_tree_0__3__8_), .A1(n26156), 
        .B0(M2_U4_U1_enc_tree_0__3__24_), .Y(M2_U4_U1_enc_tree_0__4__16_) );
  OAI21XL M2_U4_U1_UEN1_0_2_3 ( .A0(M2_U4_U1_enc_tree_0__1__26_), .A1(
        M2_U4_U1_or2_inv_0__28_), .B0(M2_U4_U1_enc_tree_0__1__30_), .Y(
        M2_U4_U1_enc_tree_0__2__28_) );
  OAI21XL M2_U4_U1_UEN1_0_2_2 ( .A0(M2_U4_U1_enc_tree_0__1__18_), .A1(
        M2_U4_U1_or2_inv_0__20_), .B0(M2_U4_U1_enc_tree_0__1__22_), .Y(
        M2_U4_U1_enc_tree_0__2__20_) );
  OAI21XL M2_U4_U1_UEN1_0_2_1 ( .A0(M2_U4_U1_enc_tree_0__1__10_), .A1(n6206), 
        .B0(M2_U4_U1_enc_tree_0__1__14_), .Y(M2_U4_U1_enc_tree_0__2__12_) );
  OAI21XL M0_U4_U1_UEN1_2_4_0 ( .A0(n25988), .A1(n26198), .B0(
        M0_U4_U1_enc_tree_2__3__24_), .Y(M0_U4_U1_enc_tree_2__4__16_) );
  OAI21XL M0_U4_U1_UEN1_1_4_0 ( .A0(M0_U4_U1_enc_tree_1__3__8_), .A1(n26148), 
        .B0(M0_U4_U1_enc_tree_1__3__24_), .Y(M0_U4_U1_enc_tree_1__4__16_) );
  OAI21XL M0_U4_U1_UEN1_1_2_3 ( .A0(M0_U4_U1_enc_tree_1__1__26_), .A1(n5576), 
        .B0(M0_U4_U1_enc_tree_1__1__30_), .Y(M0_U4_U1_enc_tree_1__2__28_) );
  OAI21XL M0_U4_U1_UEN1_1_2_2 ( .A0(M0_U4_U1_enc_tree_1__1__18_), .A1(
        M0_U4_U1_or2_inv_1__20_), .B0(M0_U4_U1_enc_tree_1__1__22_), .Y(
        M0_U4_U1_enc_tree_1__2__20_) );
  OAI21XL M0_U4_U1_UEN1_1_2_1 ( .A0(M0_U4_U1_enc_tree_1__1__10_), .A1(
        M0_U4_U1_or2_inv_1__12_), .B0(M0_U4_U1_enc_tree_1__1__14_), .Y(
        M0_U4_U1_enc_tree_1__2__12_) );
  OAI21XL M0_U4_U1_UEN1_0_4_0 ( .A0(M0_U4_U1_enc_tree_0__3__8_), .A1(n26149), 
        .B0(M0_U4_U1_enc_tree_0__3__24_), .Y(M0_U4_U1_enc_tree_0__4__16_) );
  OAI21XL M0_U4_U1_UEN1_0_2_3 ( .A0(M0_U4_U1_enc_tree_0__1__26_), .A1(n5577), 
        .B0(M0_U4_U1_enc_tree_0__1__30_), .Y(M0_U4_U1_enc_tree_0__2__28_) );
  OAI21XL M0_U4_U1_UEN1_0_2_2 ( .A0(M0_U4_U1_enc_tree_0__1__18_), .A1(
        M0_U4_U1_or2_inv_0__20_), .B0(M0_U4_U1_enc_tree_0__1__22_), .Y(
        M0_U4_U1_enc_tree_0__2__20_) );
  OAI21XL M0_U4_U1_UEN1_0_2_1 ( .A0(M0_U4_U1_enc_tree_0__1__10_), .A1(
        M0_U4_U1_or2_tree_0__1__12_), .B0(M0_U4_U1_enc_tree_0__1__14_), .Y(
        M0_U4_U1_enc_tree_0__2__12_) );
  OAI21XL M1_U4_U1_UEN1_2_4_0 ( .A0(n25983), .A1(n26202), .B0(
        M1_U4_U1_enc_tree_2__3__24_), .Y(M1_U4_U1_enc_tree_2__4__16_) );
  OAI21XL M1_U4_U1_UEN1_1_4_0 ( .A0(M1_U4_U1_enc_tree_1__3__8_), .A1(n26211), 
        .B0(M1_U4_U1_enc_tree_1__3__24_), .Y(M1_U4_U1_enc_tree_1__4__16_) );
  OAI21XL M1_U4_U1_UEN1_1_2_3 ( .A0(M1_U4_U1_enc_tree_1__1__26_), .A1(
        M1_U4_U1_or2_inv_1__28_), .B0(M1_U4_U1_enc_tree_1__1__30_), .Y(
        M1_U4_U1_enc_tree_1__2__28_) );
  OAI21XL M1_U4_U1_UEN1_1_2_2 ( .A0(M1_U4_U1_enc_tree_1__1__18_), .A1(
        M1_U4_U1_or2_inv_1__20_), .B0(M1_U4_U1_enc_tree_1__1__22_), .Y(
        M1_U4_U1_enc_tree_1__2__20_) );
  OAI21XL M1_U4_U1_UEN1_1_2_1 ( .A0(M1_U4_U1_enc_tree_1__1__10_), .A1(
        M1_U4_U1_or2_inv_1__12_), .B0(M1_U4_U1_enc_tree_1__1__14_), .Y(
        M1_U4_U1_enc_tree_1__2__12_) );
  OAI21XL M1_U4_U1_UEN1_0_4_0 ( .A0(M1_U4_U1_enc_tree_0__3__8_), .A1(n26212), 
        .B0(M1_U4_U1_enc_tree_0__3__24_), .Y(M1_U4_U1_enc_tree_0__4__16_) );
  OAI21XL M1_U4_U1_UEN1_0_2_3 ( .A0(M1_U4_U1_enc_tree_0__1__26_), .A1(
        M1_U4_U1_or2_inv_0__28_), .B0(M1_U4_U1_enc_tree_0__1__30_), .Y(
        M1_U4_U1_enc_tree_0__2__28_) );
  OAI21XL M1_U4_U1_UEN1_0_2_2 ( .A0(M1_U4_U1_enc_tree_0__1__18_), .A1(
        M1_U4_U1_or2_inv_0__20_), .B0(M1_U4_U1_enc_tree_0__1__22_), .Y(
        M1_U4_U1_enc_tree_0__2__20_) );
  OAI21XL M1_U4_U1_UEN1_0_2_1 ( .A0(M1_U4_U1_enc_tree_0__1__10_), .A1(
        M1_U4_U1_or2_tree_0__1__12_), .B0(M1_U4_U1_enc_tree_0__1__14_), .Y(
        M1_U4_U1_enc_tree_0__2__12_) );
  AOI21XL M1_U4_U1_UEN0_0_1_7 ( .A0(M1_b_2_), .A1(n3214), .B0(M1_b_0_), .Y(
        M1_U4_U1_enc_tree_0__1__30_) );
  AOI21XL M1_U4_U1_UEN0_0_1_2 ( .A0(M1_b_22_), .A1(n14290), .B0(M1_b_20_), .Y(
        M1_U4_U1_enc_tree_0__1__10_) );
  OAI21XL M0_U3_U1_UEN1_2_4_0 ( .A0(n25986), .A1(n26201), .B0(
        M0_U3_U1_enc_tree_2__3__24_), .Y(M0_U3_U1_enc_tree_2__4__16_) );
  OAI21XL M0_U3_U1_UEN1_1_4_0 ( .A0(M0_U3_U1_enc_tree_1__3__8_), .A1(n26147), 
        .B0(M0_U3_U1_enc_tree_1__3__24_), .Y(M0_U3_U1_enc_tree_1__4__16_) );
  OAI21XL M0_U3_U1_UEN1_1_2_3 ( .A0(M0_U3_U1_enc_tree_1__1__26_), .A1(
        M0_U3_U1_or2_inv_1__28_), .B0(M0_U3_U1_enc_tree_1__1__30_), .Y(
        M0_U3_U1_enc_tree_1__2__28_) );
  OAI21XL M0_U3_U1_UEN1_1_2_2 ( .A0(M0_U3_U1_enc_tree_1__1__18_), .A1(
        M0_U3_U1_or2_inv_1__20_), .B0(M0_U3_U1_enc_tree_1__1__22_), .Y(
        M0_U3_U1_enc_tree_1__2__20_) );
  OAI21XL M0_U3_U1_UEN1_1_2_1 ( .A0(M0_U3_U1_enc_tree_1__1__10_), .A1(
        M0_U3_U1_or2_inv_1__12_), .B0(M0_U3_U1_enc_tree_1__1__14_), .Y(
        M0_U3_U1_enc_tree_1__2__12_) );
  OAI21XL M0_U3_U1_UEN1_0_4_0 ( .A0(M0_U3_U1_enc_tree_0__3__8_), .A1(n26152), 
        .B0(M0_U3_U1_enc_tree_0__3__24_), .Y(M0_U3_U1_enc_tree_0__4__16_) );
  OAI21XL M0_U3_U1_UEN1_0_2_3 ( .A0(M0_U3_U1_enc_tree_0__1__26_), .A1(
        M0_U3_U1_or2_inv_0__28_), .B0(M0_U3_U1_enc_tree_0__1__30_), .Y(
        M0_U3_U1_enc_tree_0__2__28_) );
  OAI21XL M0_U3_U1_UEN1_0_2_2 ( .A0(M0_U3_U1_enc_tree_0__1__18_), .A1(
        M0_U3_U1_or2_inv_0__20_), .B0(M0_U3_U1_enc_tree_0__1__22_), .Y(
        M0_U3_U1_enc_tree_0__2__20_) );
  OAI21XL M0_U3_U1_UEN1_0_2_1 ( .A0(M0_U3_U1_enc_tree_0__1__10_), .A1(
        M0_U3_U1_or2_tree_0__1__12_), .B0(M0_U3_U1_enc_tree_0__1__14_), .Y(
        M0_U3_U1_enc_tree_0__2__12_) );
  OAI21XL M4_U3_U1_UEN1_2_4_0 ( .A0(n25985), .A1(n26200), .B0(
        M4_U3_U1_enc_tree_2__3__24_), .Y(M4_U3_U1_enc_tree_2__4__16_) );
  OAI21XL M4_U3_U1_UEN1_1_4_0 ( .A0(M4_U3_U1_enc_tree_1__3__8_), .A1(n26150), 
        .B0(M4_U3_U1_enc_tree_1__3__24_), .Y(M4_U3_U1_enc_tree_1__4__16_) );
  OAI21XL M4_U3_U1_UEN1_1_2_3 ( .A0(M4_U3_U1_enc_tree_1__1__26_), .A1(
        M4_U3_U1_or2_inv_1__28_), .B0(M4_U3_U1_enc_tree_1__1__30_), .Y(
        M4_U3_U1_enc_tree_1__2__28_) );
  OAI21XL M4_U3_U1_UEN1_1_2_2 ( .A0(M4_U3_U1_enc_tree_1__1__18_), .A1(
        M4_U3_U1_or2_inv_1__20_), .B0(M4_U3_U1_enc_tree_1__1__22_), .Y(
        M4_U3_U1_enc_tree_1__2__20_) );
  OAI21XL M4_U3_U1_UEN1_1_2_1 ( .A0(M4_U3_U1_enc_tree_1__1__10_), .A1(
        M4_U3_U1_or2_inv_1__12_), .B0(M4_U3_U1_enc_tree_1__1__14_), .Y(
        M4_U3_U1_enc_tree_1__2__12_) );
  OAI21XL M4_U3_U1_UEN1_0_4_0 ( .A0(M4_U3_U1_enc_tree_0__3__8_), .A1(n26154), 
        .B0(M4_U3_U1_enc_tree_0__3__24_), .Y(M4_U3_U1_enc_tree_0__4__16_) );
  OAI21XL M4_U3_U1_UEN1_0_2_3 ( .A0(M4_U3_U1_enc_tree_0__1__26_), .A1(
        M4_U3_U1_or2_inv_0__28_), .B0(M4_U3_U1_enc_tree_0__1__30_), .Y(
        M4_U3_U1_enc_tree_0__2__28_) );
  OAI21XL M4_U3_U1_UEN1_0_2_2 ( .A0(M4_U3_U1_enc_tree_0__1__18_), .A1(
        M4_U3_U1_or2_inv_0__20_), .B0(M4_U3_U1_enc_tree_0__1__22_), .Y(
        M4_U3_U1_enc_tree_0__2__20_) );
  OAI21XL M4_U3_U1_UEN1_0_2_1 ( .A0(M4_U3_U1_enc_tree_0__1__10_), .A1(
        M4_U3_U1_or2_tree_0__1__12_), .B0(M4_U3_U1_enc_tree_0__1__14_), .Y(
        M4_U3_U1_enc_tree_0__2__12_) );
  OAI21XL M3_U3_U1_UEN1_2_4_0 ( .A0(n25990), .A1(n26203), .B0(
        M3_U3_U1_enc_tree_2__3__24_), .Y(M3_U3_U1_enc_tree_2__4__16_) );
  OAI21XL M3_U3_U1_UEN1_1_4_0 ( .A0(M3_U3_U1_enc_tree_1__3__8_), .A1(n26151), 
        .B0(M3_U3_U1_enc_tree_1__3__24_), .Y(M3_U3_U1_enc_tree_1__4__16_) );
  OAI21XL M3_U3_U1_UEN1_1_2_3 ( .A0(M3_U3_U1_enc_tree_1__1__26_), .A1(
        M3_U3_U1_or2_inv_1__28_), .B0(M3_U3_U1_enc_tree_1__1__30_), .Y(
        M3_U3_U1_enc_tree_1__2__28_) );
  OAI21XL M3_U3_U1_UEN1_1_2_2 ( .A0(M3_U3_U1_enc_tree_1__1__18_), .A1(
        M3_U3_U1_or2_inv_1__20_), .B0(M3_U3_U1_enc_tree_1__1__22_), .Y(
        M3_U3_U1_enc_tree_1__2__20_) );
  OAI21XL M3_U3_U1_UEN1_1_2_1 ( .A0(M3_U3_U1_enc_tree_1__1__10_), .A1(
        M3_U3_U1_or2_inv_1__12_), .B0(M3_U3_U1_enc_tree_1__1__14_), .Y(
        M3_U3_U1_enc_tree_1__2__12_) );
  OAI21XL M3_U3_U1_UEN1_0_4_0 ( .A0(M3_U3_U1_enc_tree_0__3__8_), .A1(n26158), 
        .B0(M3_U3_U1_enc_tree_0__3__24_), .Y(M3_U3_U1_enc_tree_0__4__16_) );
  OAI21XL M3_U3_U1_UEN1_0_2_3 ( .A0(M3_U3_U1_enc_tree_0__1__26_), .A1(
        M3_U3_U1_or2_inv_0__28_), .B0(M3_U3_U1_enc_tree_0__1__30_), .Y(
        M3_U3_U1_enc_tree_0__2__28_) );
  OAI21XL M3_U3_U1_UEN1_0_2_2 ( .A0(M3_U3_U1_enc_tree_0__1__18_), .A1(
        M3_U3_U1_or2_inv_0__20_), .B0(M3_U3_U1_enc_tree_0__1__22_), .Y(
        M3_U3_U1_enc_tree_0__2__20_) );
  OAI21XL M3_U3_U1_UEN1_0_2_1 ( .A0(M3_U3_U1_enc_tree_0__1__10_), .A1(n4693), 
        .B0(M3_U3_U1_enc_tree_0__1__14_), .Y(M3_U3_U1_enc_tree_0__2__12_) );
  OAI21XL M5_U3_U1_UEN1_2_4_0 ( .A0(n25982), .A1(n26196), .B0(
        M5_U3_U1_enc_tree_2__3__24_), .Y(M5_U3_U1_enc_tree_2__4__16_) );
  OAI21XL M5_U3_U1_UEN1_1_4_0 ( .A0(M5_U3_U1_enc_tree_1__3__8_), .A1(n26206), 
        .B0(M5_U3_U1_enc_tree_1__3__24_), .Y(M5_U3_U1_enc_tree_1__4__16_) );
  OAI21XL M5_U3_U1_UEN1_1_2_3 ( .A0(M5_U3_U1_enc_tree_1__1__26_), .A1(
        M5_U3_U1_or2_inv_1__28_), .B0(M5_U3_U1_enc_tree_1__1__30_), .Y(
        M5_U3_U1_enc_tree_1__2__28_) );
  OAI21XL M5_U3_U1_UEN1_1_2_2 ( .A0(M5_U3_U1_enc_tree_1__1__18_), .A1(
        M5_U3_U1_or2_inv_1__20_), .B0(M5_U3_U1_enc_tree_1__1__22_), .Y(
        M5_U3_U1_enc_tree_1__2__20_) );
  OAI21XL M5_U3_U1_UEN1_1_2_1 ( .A0(M5_U3_U1_enc_tree_1__1__10_), .A1(
        M5_U3_U1_or2_inv_1__12_), .B0(M5_U3_U1_enc_tree_1__1__14_), .Y(
        M5_U3_U1_enc_tree_1__2__12_) );
  OAI21XL M5_U3_U1_UEN1_0_4_0 ( .A0(M5_U3_U1_enc_tree_0__3__8_), .A1(n26208), 
        .B0(M5_U3_U1_enc_tree_0__3__24_), .Y(M5_U3_U1_enc_tree_0__4__16_) );
  OAI21XL M5_U3_U1_UEN1_0_2_3 ( .A0(M5_U3_U1_enc_tree_0__1__26_), .A1(
        M5_U3_U1_or2_inv_0__28_), .B0(M5_U3_U1_enc_tree_0__1__30_), .Y(
        M5_U3_U1_enc_tree_0__2__28_) );
  OAI21XL M5_U3_U1_UEN1_0_2_2 ( .A0(M5_U3_U1_enc_tree_0__1__18_), .A1(
        M5_U3_U1_or2_inv_0__20_), .B0(M5_U3_U1_enc_tree_0__1__22_), .Y(
        M5_U3_U1_enc_tree_0__2__20_) );
  OAI21XL M5_U3_U1_UEN1_0_2_1 ( .A0(M5_U3_U1_enc_tree_0__1__10_), .A1(n4694), 
        .B0(M5_U3_U1_enc_tree_0__1__14_), .Y(M5_U3_U1_enc_tree_0__2__12_) );
  OAI21XL M4_U4_U1_UEN1_1_2_1 ( .A0(M4_U4_U1_enc_tree_1__1__10_), .A1(
        M4_U4_U1_or2_inv_1__12_), .B0(M4_U4_U1_enc_tree_1__1__14_), .Y(
        M4_U4_U1_enc_tree_1__2__12_) );
  OAI21XL M4_U4_U1_UEN1_0_2_1 ( .A0(M4_U4_U1_enc_tree_0__1__10_), .A1(
        M4_U4_U1_or2_tree_0__1__12_), .B0(M4_U4_U1_enc_tree_0__1__14_), .Y(
        M4_U4_U1_enc_tree_0__2__12_) );
  AOI21XL M4_U4_U1_UEN0_0_1_3 ( .A0(n3196), .A1(M4_U4_U1_or2_inv_0__14_), .B0(
        n11495), .Y(M4_U4_U1_enc_tree_0__1__14_) );
  OAI21XL M3_U4_U1_UEN1_2_4_0 ( .A0(n25893), .A1(n26146), .B0(
        M3_U4_U1_enc_tree_2__3__24_), .Y(M3_U4_U1_enc_tree_2__4__16_) );
  OAI21XL M3_U4_U1_UEN1_1_4_0 ( .A0(M3_U4_U1_enc_tree_1__3__8_), .A1(n26155), 
        .B0(M3_U4_U1_enc_tree_1__3__24_), .Y(M3_U4_U1_enc_tree_1__4__16_) );
  OAI21XL M3_U4_U1_UEN1_1_2_3 ( .A0(M4_U4_U1_enc_tree_1__1__26_), .A1(
        M3_U4_U1_or2_inv_1__28_), .B0(M4_U4_U1_enc_tree_1__1__30_), .Y(
        M3_U4_U1_enc_tree_1__2__28_) );
  OAI21XL M3_U4_U1_UEN1_1_2_2 ( .A0(M4_U4_U1_enc_tree_1__1__18_), .A1(
        M3_U4_U1_or2_inv_1__20_), .B0(M4_U4_U1_enc_tree_1__1__22_), .Y(
        M3_U4_U1_enc_tree_1__2__20_) );
  OAI21XL M3_U4_U1_UEN1_0_4_0 ( .A0(M3_U4_U1_enc_tree_0__3__8_), .A1(n26157), 
        .B0(M3_U4_U1_enc_tree_0__3__24_), .Y(M3_U4_U1_enc_tree_0__4__16_) );
  OAI21XL M3_U4_U1_UEN1_0_2_3 ( .A0(M3_U4_U1_enc_tree_0__1__26_), .A1(
        M3_U4_U1_or2_inv_0__28_), .B0(M3_U4_U1_enc_tree_0__1__30_), .Y(
        M3_U4_U1_enc_tree_0__2__28_) );
  OAI21XL M3_U4_U1_UEN1_0_2_2 ( .A0(M3_U4_U1_enc_tree_0__1__18_), .A1(
        M3_U4_U1_or2_inv_0__20_), .B0(M3_U4_U1_enc_tree_0__1__22_), .Y(
        M3_U4_U1_enc_tree_0__2__20_) );
  DFFSX1 w1_reg_11__30_ ( .D(n2130), .CK(clk), .SN(rst_n), .Q(n26485), .QN(
        w1[382]) );
  DFFSX1 w1_reg_11__29_ ( .D(n2126), .CK(clk), .SN(rst_n), .Q(n26460), .QN(
        w1[381]) );
  DFFSX1 w1_reg_11__26_ ( .D(n2114), .CK(clk), .SN(rst_n), .Q(n26457), .QN(
        w1[378]) );
  DFFSX1 w1_reg_11__25_ ( .D(n2110), .CK(clk), .SN(rst_n), .Q(n26459), .QN(
        w1[377]) );
  DFFSX1 w1_reg_11__24_ ( .D(n2106), .CK(clk), .SN(rst_n), .Q(n26461), .QN(
        w1[376]) );
  DFFSX1 w1_reg_11__23_ ( .D(n2102), .CK(clk), .SN(rst_n), .Q(n26458), .QN(
        w1[375]) );
  DFFSX1 w1_reg_11__22_ ( .D(n2098), .CK(clk), .SN(rst_n), .Q(n26462), .QN(
        w1[374]) );
  DFFSX1 w1_reg_11__21_ ( .D(n2094), .CK(clk), .SN(rst_n), .Q(n26463), .QN(
        w1[373]) );
  DFFSX1 w1_reg_11__20_ ( .D(n2090), .CK(clk), .SN(rst_n), .Q(n26464), .QN(
        w1[372]) );
  DFFSX1 w1_reg_11__19_ ( .D(n2086), .CK(clk), .SN(rst_n), .Q(n26465), .QN(
        w1[371]) );
  DFFSX1 w1_reg_11__18_ ( .D(n2082), .CK(clk), .SN(rst_n), .Q(n26466), .QN(
        w1[370]) );
  DFFSX1 w1_reg_11__17_ ( .D(n2078), .CK(clk), .SN(rst_n), .Q(n26467), .QN(
        w1[369]) );
  DFFSX1 w1_reg_11__16_ ( .D(n2074), .CK(clk), .SN(rst_n), .Q(n26468), .QN(
        w1[368]) );
  DFFSX1 w1_reg_11__15_ ( .D(n2070), .CK(clk), .SN(rst_n), .Q(n26469), .QN(
        w1[367]) );
  DFFSX1 w1_reg_11__14_ ( .D(n2066), .CK(clk), .SN(rst_n), .Q(n26470), .QN(
        w1[366]) );
  DFFSX1 w1_reg_11__13_ ( .D(n2062), .CK(clk), .SN(rst_n), .Q(n26471), .QN(
        w1[365]) );
  DFFSX1 w1_reg_11__12_ ( .D(n2058), .CK(clk), .SN(rst_n), .Q(n26472), .QN(
        w1[364]) );
  DFFSX1 w1_reg_11__11_ ( .D(n2054), .CK(clk), .SN(rst_n), .Q(n26473), .QN(
        w1[363]) );
  DFFSX1 w1_reg_11__10_ ( .D(n2050), .CK(clk), .SN(rst_n), .Q(n26474), .QN(
        w1[362]) );
  DFFSX1 w1_reg_11__9_ ( .D(n2046), .CK(clk), .SN(rst_n), .Q(n26475), .QN(
        w1[361]) );
  DFFSX1 w1_reg_11__8_ ( .D(n2042), .CK(clk), .SN(rst_n), .Q(n26476), .QN(
        w1[360]) );
  DFFSX1 w1_reg_11__7_ ( .D(n2038), .CK(clk), .SN(rst_n), .Q(n26477), .QN(
        w1[359]) );
  DFFSX1 w1_reg_11__6_ ( .D(n2034), .CK(clk), .SN(rst_n), .Q(n26478), .QN(
        w1[358]) );
  DFFSX1 w1_reg_11__5_ ( .D(n2030), .CK(clk), .SN(rst_n), .Q(n26479), .QN(
        w1[357]) );
  DFFSX1 w1_reg_11__4_ ( .D(n2026), .CK(clk), .SN(rst_n), .Q(n26480), .QN(
        w1[356]) );
  DFFSX1 w1_reg_11__3_ ( .D(n2022), .CK(clk), .SN(rst_n), .Q(n26481), .QN(
        w1[355]) );
  DFFSX1 w1_reg_11__2_ ( .D(n2018), .CK(clk), .SN(rst_n), .Q(n26482), .QN(
        w1[354]) );
  DFFSX1 w1_reg_11__1_ ( .D(n2014), .CK(clk), .SN(rst_n), .Q(n26483), .QN(
        w1[353]) );
  DFFSX1 w1_reg_11__0_ ( .D(n2010), .CK(clk), .SN(rst_n), .Q(n26484), .QN(
        w1[352]) );
  DFFSX1 w1_reg_10__22_ ( .D(n2097), .CK(clk), .SN(rst_n), .Q(n26115), .QN(
        w1[342]) );
  DFFSX1 w1_reg_10__21_ ( .D(n2093), .CK(clk), .SN(rst_n), .Q(n26116), .QN(
        w1[341]) );
  DFFSX1 w1_reg_10__20_ ( .D(n2089), .CK(clk), .SN(rst_n), .Q(n26117), .QN(
        w1[340]) );
  DFFSX1 w1_reg_10__19_ ( .D(n2085), .CK(clk), .SN(rst_n), .Q(n26118), .QN(
        w1[339]) );
  DFFSX1 w1_reg_10__18_ ( .D(n2081), .CK(clk), .SN(rst_n), .Q(n26119), .QN(
        w1[338]) );
  DFFSX1 w1_reg_10__17_ ( .D(n2077), .CK(clk), .SN(rst_n), .Q(n26120), .QN(
        w1[337]) );
  DFFSX1 w1_reg_10__15_ ( .D(n2069), .CK(clk), .SN(rst_n), .Q(n26121), .QN(
        w1[335]) );
  DFFSX1 w1_reg_10__14_ ( .D(n2065), .CK(clk), .SN(rst_n), .Q(n26122), .QN(
        w1[334]) );
  DFFSX1 w1_reg_10__13_ ( .D(n2061), .CK(clk), .SN(rst_n), .Q(n26123), .QN(
        w1[333]) );
  DFFSX1 w1_reg_10__12_ ( .D(n2057), .CK(clk), .SN(rst_n), .Q(n26136), .QN(
        w1[332]) );
  DFFSX1 w1_reg_10__11_ ( .D(n2053), .CK(clk), .SN(rst_n), .Q(n26124), .QN(
        w1[331]) );
  DFFSX1 w1_reg_10__10_ ( .D(n2049), .CK(clk), .SN(rst_n), .Q(n26125), .QN(
        w1[330]) );
  DFFSX1 w1_reg_10__3_ ( .D(n2021), .CK(clk), .SN(rst_n), .Q(n26130), .QN(
        w1[323]) );
  DFFSX1 w1_reg_10__2_ ( .D(n2017), .CK(clk), .SN(rst_n), .Q(n26131), .QN(
        w1[322]) );
  DFFSX1 w1_reg_10__1_ ( .D(n2013), .CK(clk), .SN(rst_n), .Q(n26132), .QN(
        w1[321]) );
  DFFSX1 w1_reg_10__0_ ( .D(n2009), .CK(clk), .SN(rst_n), .Q(n26133), .QN(
        w1[320]) );
  DFFSX1 w1_reg_10__9_ ( .D(n2045), .CK(clk), .SN(rst_n), .Q(n26060), .QN(
        w1[329]) );
  DFFSX1 w1_reg_10__8_ ( .D(n2041), .CK(clk), .SN(rst_n), .Q(n26061), .QN(
        w1[328]) );
  DFFSX1 w1_reg_11__28_ ( .D(n2122), .CK(clk), .SN(rst_n), .Q(n26486), .QN(
        w1[380]) );
  DFFSX1 w1_reg_11__27_ ( .D(n2118), .CK(clk), .SN(rst_n), .Q(n26413), .QN(
        w1[379]) );
  DFFSX1 w1_reg_9__9_ ( .D(n2044), .CK(clk), .SN(rst_n), .Q(n26534), .QN(
        w1[297]) );
  DFFSX1 w1_reg_9__8_ ( .D(n2040), .CK(clk), .SN(rst_n), .Q(n26536), .QN(
        w1[296]) );
  DFFSX1 w1_reg_9__22_ ( .D(n2096), .CK(clk), .SN(rst_n), .QN(w1[310]) );
  DFFSX1 w1_reg_9__29_ ( .D(n2124), .CK(clk), .SN(rst_n), .QN(w1[317]) );
  DFFSX1 w1_reg_9__28_ ( .D(n2120), .CK(clk), .SN(rst_n), .QN(w1[316]) );
  DFFSX1 w1_reg_9__24_ ( .D(n2104), .CK(clk), .SN(rst_n), .QN(w1[312]) );
  DFFSX1 w1_reg_9__23_ ( .D(n2100), .CK(clk), .SN(rst_n), .QN(w1[311]) );
  DFFSX1 w1_reg_9__21_ ( .D(n2092), .CK(clk), .SN(rst_n), .QN(w1[309]) );
  DFFSX1 w1_reg_9__20_ ( .D(n2088), .CK(clk), .SN(rst_n), .QN(w1[308]) );
  DFFSX1 w1_reg_9__19_ ( .D(n2084), .CK(clk), .SN(rst_n), .QN(w1[307]) );
  DFFSX1 w1_reg_9__17_ ( .D(n2076), .CK(clk), .SN(rst_n), .QN(w1[305]) );
  DFFSX1 w1_reg_9__16_ ( .D(n2072), .CK(clk), .SN(rst_n), .QN(w1[304]) );
  DFFSX1 w1_reg_9__15_ ( .D(n2068), .CK(clk), .SN(rst_n), .QN(w1[303]) );
  DFFSX1 w1_reg_9__14_ ( .D(n2064), .CK(clk), .SN(rst_n), .QN(w1[302]) );
  DFFSX1 w1_reg_9__11_ ( .D(n2052), .CK(clk), .SN(rst_n), .QN(w1[299]) );
  DFFSX1 w1_reg_9__10_ ( .D(n2048), .CK(clk), .SN(rst_n), .QN(w1[298]) );
  DFFSX1 w1_reg_9__7_ ( .D(n2036), .CK(clk), .SN(rst_n), .QN(w1[295]) );
  DFFSX1 w1_reg_9__6_ ( .D(n2032), .CK(clk), .SN(rst_n), .QN(w1[294]) );
  DFFSX1 w1_reg_9__5_ ( .D(n2028), .CK(clk), .SN(rst_n), .QN(w1[293]) );
  DFFSX1 w1_reg_9__4_ ( .D(n2024), .CK(clk), .SN(rst_n), .QN(w1[292]) );
  DFFSX1 w1_reg_9__3_ ( .D(n2020), .CK(clk), .SN(rst_n), .QN(w1[291]) );
  DFFSX1 w1_reg_9__1_ ( .D(n2012), .CK(clk), .SN(rst_n), .QN(w1[289]) );
  DFFSX1 w1_reg_9__12_ ( .D(n2056), .CK(clk), .SN(rst_n), .QN(w1[300]) );
  DFFSX1 w1_reg_9__30_ ( .D(n2128), .CK(clk), .SN(rst_n), .QN(w1[318]) );
  DFFSX1 w1_reg_10__27_ ( .D(n2117), .CK(clk), .SN(rst_n), .QN(w1[347]) );
  DFFSX1 w1_reg_9__27_ ( .D(n2116), .CK(clk), .SN(rst_n), .QN(w1[315]) );
  DFFSX1 w1_reg_9__26_ ( .D(n2112), .CK(clk), .SN(rst_n), .QN(w1[314]) );
  DFFSX1 w1_reg_9__25_ ( .D(n2108), .CK(clk), .SN(rst_n), .QN(w1[313]) );
  DFFSX1 w1_reg_9__18_ ( .D(n2080), .CK(clk), .SN(rst_n), .QN(w1[306]) );
  DFFSX1 w1_reg_9__13_ ( .D(n2060), .CK(clk), .SN(rst_n), .QN(w1[301]) );
  DFFSX1 w1_reg_9__2_ ( .D(n2016), .CK(clk), .SN(rst_n), .QN(w1[290]) );
  DFFSX1 w1_reg_9__0_ ( .D(n2008), .CK(clk), .SN(rst_n), .QN(w1[288]) );
  DFFSX1 sigma11_reg_30_ ( .D(n2357), .CK(clk), .SN(rst_n), .Q(n26108), .QN(
        sigma11[30]) );
  DFFSX1 sigma11_reg_29_ ( .D(n2355), .CK(clk), .SN(rst_n), .Q(n26139), .QN(
        sigma11[29]) );
  DFFSX1 sigma11_reg_28_ ( .D(n2353), .CK(clk), .SN(rst_n), .Q(n26106), .QN(
        sigma11[28]) );
  DFFSX1 sigma11_reg_27_ ( .D(n2351), .CK(clk), .SN(rst_n), .Q(n26455), .QN(
        sigma11[27]) );
  DFFSX1 sigma12_reg_30_ ( .D(n2356), .CK(clk), .SN(rst_n), .Q(n26454), .QN(
        sigma12[30]) );
  DFFSX1 sigma12_reg_28_ ( .D(n2352), .CK(clk), .SN(rst_n), .Q(n26452), .QN(
        sigma12[28]) );
  DFFSX1 sigma12_reg_27_ ( .D(n2350), .CK(clk), .SN(rst_n), .Q(n26519), .QN(
        sigma12[27]) );
  DFFSX1 sigma11_reg_26_ ( .D(n2349), .CK(clk), .SN(rst_n), .Q(n26456), .QN(
        sigma11[26]) );
  DFFSX1 sigma11_reg_25_ ( .D(n2347), .CK(clk), .SN(rst_n), .Q(n26138), .QN(
        sigma11[25]) );
  DFFSX1 sigma12_reg_26_ ( .D(n2348), .CK(clk), .SN(rst_n), .Q(n6220), .QN(
        sigma12[26]) );
  DFFSX1 sigma12_reg_4_ ( .D(n2304), .CK(clk), .SN(rst_n), .Q(n26041), .QN(
        sigma12[4]) );
  DFFSX1 sigma12_reg_12_ ( .D(n2320), .CK(clk), .SN(rst_n), .Q(n26518), .QN(
        sigma12[12]) );
  DFFSX1 sigma12_reg_10_ ( .D(n2316), .CK(clk), .SN(rst_n), .Q(n26516), .QN(
        sigma12[10]) );
  DFFSX1 sigma11_reg_24_ ( .D(n2345), .CK(clk), .SN(rst_n), .Q(n26416), .QN(
        sigma11[24]) );
  DFFSX1 sigma11_reg_23_ ( .D(n2343), .CK(clk), .SN(rst_n), .Q(n26107), .QN(
        sigma11[23]) );
  DFFSX1 sigma11_reg_22_ ( .D(n2341), .CK(clk), .SN(rst_n), .Q(n26451), .QN(
        sigma11[22]) );
  DFFSX1 sigma11_reg_4_ ( .D(n2305), .CK(clk), .SN(rst_n), .Q(n26370), .QN(
        sigma11[4]) );
  DFFSX1 sigma12_reg_13_ ( .D(n2322), .CK(clk), .SN(rst_n), .Q(n26032), .QN(
        sigma12[13]) );
  DFFSX1 sigma12_reg_0_ ( .D(n2296), .CK(clk), .SN(rst_n), .Q(n26513), .QN(
        sigma12[0]) );
  DFFSX1 sigma11_reg_20_ ( .D(n2337), .CK(clk), .SN(rst_n), .QN(sigma11[20])
         );
  DFFSX1 sigma11_reg_2_ ( .D(n2301), .CK(clk), .SN(rst_n), .QN(sigma11[2]) );
  DFFSX1 sigma11_reg_19_ ( .D(n2335), .CK(clk), .SN(rst_n), .QN(sigma11[19])
         );
  DFFSX1 sigma11_reg_3_ ( .D(n2303), .CK(clk), .SN(rst_n), .QN(sigma11[3]) );
  DFFSX1 out_reg_31_ ( .D(n2492), .CK(clk), .SN(rst_n), .QN(out[31]) );
  DFFSX1 out_reg_30_ ( .D(n2493), .CK(clk), .SN(rst_n), .QN(out[30]) );
  DFFSX1 out_reg_29_ ( .D(n2494), .CK(clk), .SN(rst_n), .QN(out[29]) );
  DFFSX1 out_reg_28_ ( .D(n2495), .CK(clk), .SN(rst_n), .QN(out[28]) );
  DFFSX1 out_reg_27_ ( .D(n2496), .CK(clk), .SN(rst_n), .QN(out[27]) );
  DFFSX1 out_reg_26_ ( .D(n2497), .CK(clk), .SN(rst_n), .QN(out[26]) );
  DFFSX1 out_reg_25_ ( .D(n2498), .CK(clk), .SN(rst_n), .QN(out[25]) );
  DFFSX1 out_reg_24_ ( .D(n2499), .CK(clk), .SN(rst_n), .QN(out[24]) );
  DFFSX1 out_reg_23_ ( .D(n2500), .CK(clk), .SN(rst_n), .QN(out[23]) );
  DFFSX1 out_reg_22_ ( .D(n2501), .CK(clk), .SN(rst_n), .QN(out[22]) );
  DFFSX1 out_reg_21_ ( .D(n2502), .CK(clk), .SN(rst_n), .QN(out[21]) );
  DFFSX1 out_reg_20_ ( .D(n2503), .CK(clk), .SN(rst_n), .QN(out[20]) );
  DFFSX1 out_reg_19_ ( .D(n2504), .CK(clk), .SN(rst_n), .QN(out[19]) );
  DFFSX1 out_reg_18_ ( .D(n2505), .CK(clk), .SN(rst_n), .QN(out[18]) );
  DFFSX1 out_reg_17_ ( .D(n2506), .CK(clk), .SN(rst_n), .QN(out[17]) );
  DFFSX1 out_reg_16_ ( .D(n2507), .CK(clk), .SN(rst_n), .QN(out[16]) );
  DFFSX1 out_reg_15_ ( .D(n2508), .CK(clk), .SN(rst_n), .QN(out[15]) );
  DFFSX1 out_reg_14_ ( .D(n2509), .CK(clk), .SN(rst_n), .QN(out[14]) );
  DFFSX1 out_reg_13_ ( .D(n2510), .CK(clk), .SN(rst_n), .QN(out[13]) );
  DFFSX1 out_reg_12_ ( .D(n2511), .CK(clk), .SN(rst_n), .QN(out[12]) );
  DFFSX1 out_reg_11_ ( .D(n2512), .CK(clk), .SN(rst_n), .QN(out[11]) );
  DFFSX1 out_reg_10_ ( .D(n2513), .CK(clk), .SN(rst_n), .QN(out[10]) );
  DFFSX1 out_reg_9_ ( .D(n2514), .CK(clk), .SN(rst_n), .QN(out[9]) );
  DFFSX1 out_reg_8_ ( .D(n2515), .CK(clk), .SN(rst_n), .QN(out[8]) );
  DFFSX1 out_reg_7_ ( .D(n2516), .CK(clk), .SN(rst_n), .QN(out[7]) );
  DFFSX1 out_reg_6_ ( .D(n2517), .CK(clk), .SN(rst_n), .QN(out[6]) );
  DFFSX1 out_reg_5_ ( .D(n2518), .CK(clk), .SN(rst_n), .QN(out[5]) );
  DFFSX1 out_reg_4_ ( .D(n2519), .CK(clk), .SN(rst_n), .QN(out[4]) );
  DFFSX1 out_reg_3_ ( .D(n2520), .CK(clk), .SN(rst_n), .QN(out[3]) );
  DFFSX1 out_reg_2_ ( .D(n2521), .CK(clk), .SN(rst_n), .QN(out[2]) );
  DFFSX1 out_reg_1_ ( .D(n2522), .CK(clk), .SN(rst_n), .QN(out[1]) );
  DFFSX1 out_reg_0_ ( .D(n2523), .CK(clk), .SN(rst_n), .QN(out[0]) );
  DFFSX1 out_valid_reg ( .D(n26487), .CK(clk), .SN(rst_n), .QN(out_valid) );
  DFFSX1 sigma12_reg_14_ ( .D(n2324), .CK(clk), .SN(rst_n), .Q(n26296), .QN(
        sigma12[14]) );
  DFFSX1 sigma12_reg_6_ ( .D(n2308), .CK(clk), .SN(rst_n), .Q(n26294), .QN(
        sigma12[6]) );
  DFFSX1 sigma12_reg_3_ ( .D(n2302), .CK(clk), .SN(rst_n), .Q(n26276), .QN(
        sigma12[3]) );
  DFFSX1 sigma12_reg_2_ ( .D(n2300), .CK(clk), .SN(rst_n), .Q(n26295), .QN(
        sigma12[2]) );
  DFFSX1 sigma12_reg_1_ ( .D(n2298), .CK(clk), .SN(rst_n), .Q(n26270), .QN(
        sigma12[1]) );
  DFFSX1 sigma12_reg_8_ ( .D(n2312), .CK(clk), .SN(rst_n), .Q(n25932), .QN(
        sigma12[8]) );
  DFFSX1 sigma12_reg_5_ ( .D(n2306), .CK(clk), .SN(rst_n), .Q(n26031), .QN(
        sigma12[5]) );
  DFFSX1 sigma10_reg_9_ ( .D(n2273), .CK(clk), .SN(rst_n), .Q(n26232), .QN(
        sigma10[9]) );
  DFFSX1 sigma12_reg_21_ ( .D(n2338), .CK(clk), .SN(rst_n), .QN(sigma12[21])
         );
  DFFSX1 sigma12_reg_20_ ( .D(n2336), .CK(clk), .SN(rst_n), .Q(n26038), .QN(
        sigma12[20]) );
  DFFSX1 sigma12_reg_19_ ( .D(n2334), .CK(clk), .SN(rst_n), .Q(n26020), .QN(
        sigma12[19]) );
  DFFSX1 sigma12_reg_18_ ( .D(n2332), .CK(clk), .SN(rst_n), .Q(n26275), .QN(
        sigma12[18]) );
  DFFSX1 sigma12_reg_17_ ( .D(n2330), .CK(clk), .SN(rst_n), .Q(n26019), .QN(
        sigma12[17]) );
  DFFSX1 sigma12_reg_15_ ( .D(n2326), .CK(clk), .SN(rst_n), .Q(n26018), .QN(
        sigma12[15]) );
  DFFSX1 sigma12_reg_7_ ( .D(n2310), .CK(clk), .SN(rst_n), .Q(n26277), .QN(
        sigma12[7]) );
  DFFSX1 sigma12_reg_11_ ( .D(n2318), .CK(clk), .SN(rst_n), .Q(n26517), .QN(
        sigma12[11]) );
  DFFSX1 sigma11_reg_16_ ( .D(n2329), .CK(clk), .SN(rst_n), .Q(n26449), .QN(
        sigma11[16]) );
  DFFSX1 sigma11_reg_12_ ( .D(n2321), .CK(clk), .SN(rst_n), .Q(n26448), .QN(
        sigma11[12]) );
  DFFSX1 sigma11_reg_11_ ( .D(n2319), .CK(clk), .SN(rst_n), .Q(n26447), .QN(
        sigma11[11]) );
  DFFSX1 sigma11_reg_10_ ( .D(n2317), .CK(clk), .SN(rst_n), .Q(n26446), .QN(
        sigma11[10]) );
  DFFSX1 sigma11_reg_8_ ( .D(n2313), .CK(clk), .SN(rst_n), .Q(n26445), .QN(
        sigma11[8]) );
  DFFSX1 sigma11_reg_5_ ( .D(n2307), .CK(clk), .SN(rst_n), .Q(n26444), .QN(
        sigma11[5]) );
  DFFSX1 sigma11_reg_0_ ( .D(n2297), .CK(clk), .SN(rst_n), .Q(n26450), .QN(
        sigma11[0]) );
  DFFSX1 sigma12_reg_9_ ( .D(n2314), .CK(clk), .SN(rst_n), .Q(n25925), .QN(
        sigma12[9]) );
  DFFSX1 sigma12_reg_16_ ( .D(n2328), .CK(clk), .SN(rst_n), .Q(n25917), .QN(
        sigma12[16]) );
  DFFSX1 sigma11_reg_13_ ( .D(n2323), .CK(clk), .SN(rst_n), .Q(n26443), .QN(
        sigma11[13]) );
  DFFSX1 sigma11_reg_9_ ( .D(n2315), .CK(clk), .SN(rst_n), .Q(n26369), .QN(
        sigma11[9]) );
  DFFSX1 sigma10_reg_13_ ( .D(n2277), .CK(clk), .SN(rst_n), .Q(n26235) );
  DFFSX1 sigma12_reg_22_ ( .D(n2340), .CK(clk), .SN(rst_n), .Q(n26547), .QN(
        sigma12[22]) );
  DFFSX1 sigma11_reg_18_ ( .D(n2333), .CK(clk), .SN(rst_n), .QN(sigma11[18])
         );
  DFFSX1 sigma11_reg_14_ ( .D(n2325), .CK(clk), .SN(rst_n), .QN(sigma11[14])
         );
  DFFSX1 sigma11_reg_21_ ( .D(n2339), .CK(clk), .SN(rst_n), .QN(sigma11[21])
         );
  DFFSX1 sigma11_reg_7_ ( .D(n2311), .CK(clk), .SN(rst_n), .QN(sigma11[7]) );
  DFFSX1 sigma11_reg_6_ ( .D(n2309), .CK(clk), .SN(rst_n), .QN(sigma11[6]) );
  DFFSX1 sigma11_reg_1_ ( .D(n2299), .CK(clk), .SN(rst_n), .QN(sigma11[1]) );
  DFFSX1 sigma10_reg_19_ ( .D(n2283), .CK(clk), .SN(rst_n), .Q(n25914), .QN(
        n4727) );
  DFFSX1 sigma11_reg_15_ ( .D(n2327), .CK(clk), .SN(rst_n), .Q(n4726), .QN(
        sigma11[15]) );
  DFFSX1 sigma10_reg_21_ ( .D(n2285), .CK(clk), .SN(rst_n), .Q(n25913), .QN(
        n4720) );
  DFFSX1 sigma10_reg_18_ ( .D(n2282), .CK(clk), .SN(rst_n), .Q(n25916), .QN(
        n3003) );
  DFFSX1 sigma10_reg_22_ ( .D(n2286), .CK(clk), .SN(rst_n), .Q(n25915) );
  DFFSX1 sigma11_reg_17_ ( .D(n2331), .CK(clk), .SN(rst_n), .Q(n4725), .QN(
        sigma11[17]) );
  DFFSX1 sigma10_reg_20_ ( .D(n2284), .CK(clk), .SN(rst_n), .Q(n25912), .QN(
        n4721) );
  DFFSX1 sigma10_reg_16_ ( .D(n2280), .CK(clk), .SN(rst_n), .Q(n25911) );
  DFFSX1 sigma10_reg_17_ ( .D(n2281), .CK(clk), .SN(rst_n), .Q(n25910), .QN(
        n4723) );
  DFFSX1 sigma10_reg_0_ ( .D(n2264), .CK(clk), .SN(rst_n), .Q(n25909) );
  DFFSX1 sigma10_reg_15_ ( .D(n2279), .CK(clk), .SN(rst_n), .Q(n25908), .QN(
        n4730) );
  DFFSX1 sigma10_reg_3_ ( .D(n2267), .CK(clk), .SN(rst_n), .Q(n25907), .QN(
        n4732) );
  DFFSX1 sigma10_reg_8_ ( .D(n2272), .CK(clk), .SN(rst_n), .Q(n25904), .QN(
        n4722) );
  DFFSX1 sigma10_reg_6_ ( .D(n2270), .CK(clk), .SN(rst_n), .Q(n25906), .QN(
        n4728) );
  DFFSX1 sigma10_reg_10_ ( .D(n2274), .CK(clk), .SN(rst_n), .Q(n25905), .QN(
        n4719) );
  DFFSX1 sigma10_reg_4_ ( .D(n2268), .CK(clk), .SN(rst_n), .Q(n25903), .QN(
        n4731) );
  DFFSX1 sigma10_reg_5_ ( .D(n2269), .CK(clk), .SN(rst_n), .Q(n25902), .QN(
        n4729) );
  DFFSX1 sigma10_reg_12_ ( .D(n2276), .CK(clk), .SN(rst_n), .Q(n25901), .QN(
        n4724) );
  DFFSX1 sigma10_reg_14_ ( .D(n2278), .CK(clk), .SN(rst_n), .Q(n25899), .QN(
        n4718) );
  DFFSX1 sigma10_reg_1_ ( .D(n2265), .CK(clk), .SN(rst_n), .Q(n25898) );
  DFFSX1 sigma10_reg_7_ ( .D(n2271), .CK(clk), .SN(rst_n), .Q(n25897), .QN(
        n4717) );
  DFFSX1 y11_reg_1_ ( .D(n2457), .CK(clk), .SN(rst_n), .Q(n25955), .QN(y11[1])
         );
  DFFSX1 y11_reg_0_ ( .D(n2456), .CK(clk), .SN(rst_n), .Q(n25956), .QN(y11[0])
         );
  DFFSX1 y12_reg_23_ ( .D(n2439), .CK(clk), .SN(rst_n), .Q(n26192), .QN(
        y12[23]) );
  DFFSX1 y12_reg_22_ ( .D(n2437), .CK(clk), .SN(rst_n), .Q(n25958), .QN(
        y12[22]) );
  DFFSX1 y12_reg_21_ ( .D(n2435), .CK(clk), .SN(rst_n), .Q(n25959), .QN(
        y12[21]) );
  DFFSX1 y12_reg_20_ ( .D(n2433), .CK(clk), .SN(rst_n), .Q(n25960), .QN(
        y12[20]) );
  DFFSX1 y12_reg_18_ ( .D(n2429), .CK(clk), .SN(rst_n), .Q(n25962), .QN(
        y12[18]) );
  DFFSX1 y12_reg_14_ ( .D(n2421), .CK(clk), .SN(rst_n), .Q(n25966), .QN(
        y12[14]) );
  DFFSX1 y12_reg_8_ ( .D(n2409), .CK(clk), .SN(rst_n), .Q(n25972), .QN(y12[8])
         );
  DFFSX1 y12_reg_7_ ( .D(n2407), .CK(clk), .SN(rst_n), .Q(n25973), .QN(y12[7])
         );
  DFFSX1 y12_reg_3_ ( .D(n2399), .CK(clk), .SN(rst_n), .Q(n25977), .QN(y12[3])
         );
  DFFSX1 y12_reg_0_ ( .D(n2393), .CK(clk), .SN(rst_n), .Q(n25980), .QN(y12[0])
         );
  DFFSX1 w2_reg_0__24_ ( .D(n2160), .CK(clk), .SN(rst_n), .Q(n26036), .QN(
        w2[24]) );
  DFFSX1 w2_reg_0__23_ ( .D(n2159), .CK(clk), .SN(rst_n), .Q(n26037), .QN(
        w2[23]) );
  DFFSX1 w2_reg_0__22_ ( .D(n2158), .CK(clk), .SN(rst_n), .Q(n26017), .QN(
        w2[22]) );
  DFFSX1 w2_reg_0__21_ ( .D(n2157), .CK(clk), .SN(rst_n), .Q(n26012), .QN(
        w2[21]) );
  DFFSX1 w2_reg_0__20_ ( .D(n2156), .CK(clk), .SN(rst_n), .Q(n26016), .QN(
        w2[20]) );
  DFFSX1 w2_reg_0__19_ ( .D(n2155), .CK(clk), .SN(rst_n), .Q(n26011), .QN(
        w2[19]) );
  DFFSX1 w2_reg_0__18_ ( .D(n2154), .CK(clk), .SN(rst_n), .Q(n26015), .QN(
        w2[18]) );
  DFFSX1 w2_reg_0__17_ ( .D(n2153), .CK(clk), .SN(rst_n), .Q(n26010), .QN(
        w2[17]) );
  DFFSX1 w2_reg_0__16_ ( .D(n2152), .CK(clk), .SN(rst_n), .Q(n26014), .QN(
        w2[16]) );
  DFFSX1 w2_reg_0__15_ ( .D(n2151), .CK(clk), .SN(rst_n), .Q(n26013), .QN(
        w2[15]) );
  DFFSX1 w2_reg_0__14_ ( .D(n2150), .CK(clk), .SN(rst_n), .Q(n26005), .QN(
        w2[14]) );
  DFFSX1 w2_reg_0__12_ ( .D(n2148), .CK(clk), .SN(rst_n), .Q(n26004), .QN(
        w2[12]) );
  DFFSX1 w2_reg_0__10_ ( .D(n2146), .CK(clk), .SN(rst_n), .Q(n25995), .QN(
        w2[10]) );
  DFFSX1 w2_reg_0__7_ ( .D(n2143), .CK(clk), .SN(rst_n), .Q(n25999), .QN(w2[7]) );
  DFFSX1 w2_reg_0__6_ ( .D(n2142), .CK(clk), .SN(rst_n), .Q(n26002), .QN(w2[6]) );
  DFFSX1 w2_reg_0__5_ ( .D(n2141), .CK(clk), .SN(rst_n), .Q(n25998), .QN(w2[5]) );
  DFFSX1 w2_reg_0__4_ ( .D(n2140), .CK(clk), .SN(rst_n), .Q(n26001), .QN(w2[4]) );
  DFFSX1 w2_reg_0__3_ ( .D(n2139), .CK(clk), .SN(rst_n), .Q(n26006), .QN(w2[3]) );
  DFFSX1 w2_reg_0__2_ ( .D(n2138), .CK(clk), .SN(rst_n), .Q(n26000), .QN(w2[2]) );
  DFFSX1 w2_reg_0__1_ ( .D(n2137), .CK(clk), .SN(rst_n), .Q(n25997), .QN(w2[1]) );
  DFFSX1 w2_reg_0__0_ ( .D(n2136), .CK(clk), .SN(rst_n), .Q(n26009), .QN(w2[0]) );
  DFFSX1 y11_reg_22_ ( .D(n2478), .CK(clk), .SN(rst_n), .Q(n25938), .QN(
        y11[22]) );
  DFFSX1 y11_reg_21_ ( .D(n2477), .CK(clk), .SN(rst_n), .Q(n25889), .QN(
        y11[21]) );
  DFFSX1 y11_reg_20_ ( .D(n2476), .CK(clk), .SN(rst_n), .Q(n25939), .QN(
        y11[20]) );
  DFFSX1 y11_reg_19_ ( .D(n2475), .CK(clk), .SN(rst_n), .Q(n25940), .QN(
        y11[19]) );
  DFFSX1 y11_reg_18_ ( .D(n2474), .CK(clk), .SN(rst_n), .Q(n25890), .QN(
        y11[18]) );
  DFFSX1 y11_reg_17_ ( .D(n2473), .CK(clk), .SN(rst_n), .Q(n25941), .QN(
        y11[17]) );
  DFFSX1 y11_reg_16_ ( .D(n2472), .CK(clk), .SN(rst_n), .Q(n25942), .QN(
        y11[16]) );
  DFFSX1 y11_reg_15_ ( .D(n2471), .CK(clk), .SN(rst_n), .Q(n25943), .QN(
        y11[15]) );
  DFFSX1 y11_reg_14_ ( .D(n2470), .CK(clk), .SN(rst_n), .Q(n25944), .QN(
        y11[14]) );
  DFFSX1 y11_reg_13_ ( .D(n2469), .CK(clk), .SN(rst_n), .Q(n25945), .QN(
        y11[13]) );
  DFFSX1 y11_reg_12_ ( .D(n2468), .CK(clk), .SN(rst_n), .Q(n25946), .QN(
        y11[12]) );
  DFFSX1 y11_reg_11_ ( .D(n2467), .CK(clk), .SN(rst_n), .Q(n25947), .QN(
        y11[11]) );
  DFFSX1 y11_reg_10_ ( .D(n2466), .CK(clk), .SN(rst_n), .Q(n25948), .QN(
        y11[10]) );
  DFFSX1 y11_reg_8_ ( .D(n2464), .CK(clk), .SN(rst_n), .Q(n25949), .QN(y11[8])
         );
  DFFSX1 y11_reg_7_ ( .D(n2463), .CK(clk), .SN(rst_n), .Q(n25892), .QN(y11[7])
         );
  DFFSX1 y11_reg_5_ ( .D(n2461), .CK(clk), .SN(rst_n), .Q(n25951), .QN(y11[5])
         );
  DFFSX1 y11_reg_4_ ( .D(n2460), .CK(clk), .SN(rst_n), .Q(n25952), .QN(y11[4])
         );
  DFFSX1 y11_reg_3_ ( .D(n2459), .CK(clk), .SN(rst_n), .Q(n25953), .QN(y11[3])
         );
  DFFSX1 w2_reg_0__30_ ( .D(n2166), .CK(clk), .SN(rst_n), .Q(n26046), .QN(
        w2[30]) );
  DFFSX1 w2_reg_0__29_ ( .D(n2165), .CK(clk), .SN(rst_n), .Q(n26047), .QN(
        w2[29]) );
  DFFSX1 w2_reg_0__28_ ( .D(n2164), .CK(clk), .SN(rst_n), .Q(n26301), .QN(
        w2[28]) );
  DFFSX1 w2_reg_0__27_ ( .D(n2163), .CK(clk), .SN(rst_n), .Q(n26045), .QN(
        w2[27]) );
  DFFSX1 w2_reg_0__26_ ( .D(n2162), .CK(clk), .SN(rst_n), .Q(n26043), .QN(
        w2[26]) );
  DFFSX1 w2_reg_0__25_ ( .D(n2161), .CK(clk), .SN(rst_n), .Q(n26042), .QN(
        w2[25]) );
  DFFSX1 w2_reg_0__13_ ( .D(n2149), .CK(clk), .SN(rst_n), .Q(n26026), .QN(
        w2[13]) );
  DFFSX1 w2_reg_0__9_ ( .D(n2145), .CK(clk), .SN(rst_n), .Q(n25996), .QN(w2[9]) );
  DFFSX1 y20_reg_30_ ( .D(n2390), .CK(clk), .SN(rst_n), .Q(n26159), .QN(
        y20[30]) );
  DFFSX1 y20_reg_29_ ( .D(n2389), .CK(clk), .SN(rst_n), .Q(n26164), .QN(
        y20[29]) );
  DFFSX1 y20_reg_28_ ( .D(n2388), .CK(clk), .SN(rst_n), .Q(n26163), .QN(
        y20[28]) );
  DFFSX1 y20_reg_27_ ( .D(n2387), .CK(clk), .SN(rst_n), .Q(n26161), .QN(
        y20[27]) );
  DFFSX1 y20_reg_26_ ( .D(n2386), .CK(clk), .SN(rst_n), .Q(n26165), .QN(
        y20[26]) );
  DFFSX1 y20_reg_25_ ( .D(n2385), .CK(clk), .SN(rst_n), .Q(n26162), .QN(
        y20[25]) );
  DFFSX1 y20_reg_24_ ( .D(n2384), .CK(clk), .SN(rst_n), .Q(n26160), .QN(
        y20[24]) );
  DFFSX1 y20_reg_23_ ( .D(n2383), .CK(clk), .SN(rst_n), .Q(n26166), .QN(
        y20[23]) );
  DFFSX1 y20_reg_20_ ( .D(n2380), .CK(clk), .SN(rst_n), .Q(n26168), .QN(
        y20[20]) );
  DFFSX1 y20_reg_19_ ( .D(n2379), .CK(clk), .SN(rst_n), .Q(n26170), .QN(
        y20[19]) );
  DFFSX1 y20_reg_18_ ( .D(n2378), .CK(clk), .SN(rst_n), .Q(n26171), .QN(
        y20[18]) );
  DFFSX1 y20_reg_17_ ( .D(n2377), .CK(clk), .SN(rst_n), .Q(n26172), .QN(
        y20[17]) );
  DFFSX1 y20_reg_16_ ( .D(n2376), .CK(clk), .SN(rst_n), .Q(n26173), .QN(
        y20[16]) );
  DFFSX1 y20_reg_15_ ( .D(n2375), .CK(clk), .SN(rst_n), .Q(n26174), .QN(
        y20[15]) );
  DFFSX1 y20_reg_13_ ( .D(n2373), .CK(clk), .SN(rst_n), .Q(n26176), .QN(
        y20[13]) );
  DFFSX1 y20_reg_11_ ( .D(n2371), .CK(clk), .SN(rst_n), .Q(n26178), .QN(
        y20[11]) );
  DFFSX1 y20_reg_10_ ( .D(n2370), .CK(clk), .SN(rst_n), .Q(n26179), .QN(
        y20[10]) );
  DFFSX1 y20_reg_8_ ( .D(n2368), .CK(clk), .SN(rst_n), .Q(n26180), .QN(y20[8])
         );
  DFFSX1 y20_reg_7_ ( .D(n2367), .CK(clk), .SN(rst_n), .Q(n26181), .QN(y20[7])
         );
  DFFSX1 y20_reg_6_ ( .D(n2366), .CK(clk), .SN(rst_n), .Q(n26182), .QN(y20[6])
         );
  DFFSX1 w2_reg_2__21_ ( .D(n2221), .CK(clk), .SN(rst_n), .Q(n25924), .QN(
        w2[85]) );
  DFFSX1 w2_reg_2__20_ ( .D(n2220), .CK(clk), .SN(rst_n), .Q(n25923), .QN(
        w2[84]) );
  DFFSX1 w2_reg_2__19_ ( .D(n2219), .CK(clk), .SN(rst_n), .Q(n25922), .QN(
        w2[83]) );
  DFFSX1 w2_reg_2__18_ ( .D(n2218), .CK(clk), .SN(rst_n), .Q(n26035), .QN(
        w2[82]) );
  DFFSX1 w2_reg_2__17_ ( .D(n2217), .CK(clk), .SN(rst_n), .Q(n25921), .QN(
        w2[81]) );
  DFFSX1 w2_reg_2__16_ ( .D(n2216), .CK(clk), .SN(rst_n), .Q(n26274), .QN(
        w2[80]) );
  DFFSX1 w2_reg_2__15_ ( .D(n2215), .CK(clk), .SN(rst_n), .Q(n25920), .QN(
        w2[79]) );
  DFFSX1 w2_reg_2__14_ ( .D(n2214), .CK(clk), .SN(rst_n), .Q(n25931), .QN(
        w2[78]) );
  DFFSX1 w2_reg_2__13_ ( .D(n2213), .CK(clk), .SN(rst_n), .Q(n26273), .QN(
        w2[77]) );
  DFFSX1 w2_reg_2__12_ ( .D(n2212), .CK(clk), .SN(rst_n), .Q(n26034), .QN(
        w2[76]) );
  DFFSX1 w2_reg_2__11_ ( .D(n2211), .CK(clk), .SN(rst_n), .Q(n26007), .QN(
        w2[75]) );
  DFFSX1 w2_reg_2__10_ ( .D(n2210), .CK(clk), .SN(rst_n), .Q(n26033), .QN(
        w2[74]) );
  DFFSX1 w2_reg_2__9_ ( .D(n2209), .CK(clk), .SN(rst_n), .Q(n26272), .QN(
        w2[73]) );
  DFFSX1 w2_reg_2__8_ ( .D(n2208), .CK(clk), .SN(rst_n), .Q(n26283), .QN(
        w2[72]) );
  DFFSX1 w2_reg_2__7_ ( .D(n2207), .CK(clk), .SN(rst_n), .Q(n25919), .QN(
        w2[71]) );
  DFFSX1 w2_reg_2__6_ ( .D(n2206), .CK(clk), .SN(rst_n), .Q(n26040), .QN(
        w2[70]) );
  DFFSX1 w2_reg_2__5_ ( .D(n2205), .CK(clk), .SN(rst_n), .Q(n26271), .QN(
        w2[69]) );
  DFFSX1 w2_reg_2__4_ ( .D(n2204), .CK(clk), .SN(rst_n), .Q(n26281), .QN(
        w2[68]) );
  DFFSX1 w2_reg_2__3_ ( .D(n2203), .CK(clk), .SN(rst_n), .Q(n25918), .QN(
        w2[67]) );
  DFFSX1 w2_reg_2__2_ ( .D(n2202), .CK(clk), .SN(rst_n), .Q(n25930), .QN(
        w2[66]) );
  DFFSX1 w2_reg_2__1_ ( .D(n2201), .CK(clk), .SN(rst_n), .Q(n25929), .QN(
        w2[65]) );
  DFFSX1 w2_reg_1__26_ ( .D(n2194), .CK(clk), .SN(rst_n), .Q(n26298), .QN(
        w2[58]) );
  DFFSX1 w2_reg_1__24_ ( .D(n2192), .CK(clk), .SN(rst_n), .Q(n26284), .QN(
        w2[56]) );
  DFFSX1 w2_reg_1__23_ ( .D(n2191), .CK(clk), .SN(rst_n), .Q(n26285), .QN(
        w2[55]) );
  DFFSX1 y12_reg_30_ ( .D(n2453), .CK(clk), .SN(rst_n), .Q(n25981), .QN(
        y12[30]) );
  DFFSX1 w2_reg_0__11_ ( .D(n2147), .CK(clk), .SN(rst_n), .Q(n26008), .QN(
        w2[11]) );
  DFFSX1 w2_reg_2__30_ ( .D(n2230), .CK(clk), .SN(rst_n), .Q(n26307), .QN(
        w2[94]) );
  DFFSX1 w2_reg_2__28_ ( .D(n2228), .CK(clk), .SN(rst_n), .Q(n26306), .QN(
        w2[92]) );
  DFFSX1 w2_reg_2__26_ ( .D(n2226), .CK(clk), .SN(rst_n), .Q(n26300), .QN(
        w2[90]) );
  DFFSX1 w2_reg_2__24_ ( .D(n2224), .CK(clk), .SN(rst_n), .Q(n26293), .QN(
        w2[88]) );
  DFFSX1 w2_reg_2__23_ ( .D(n2223), .CK(clk), .SN(rst_n), .Q(n26292), .QN(
        w2[87]) );
  DFFSX1 w2_reg_1__0_ ( .D(n2168), .CK(clk), .SN(rst_n), .Q(n26424), .QN(
        w2[32]) );
  DFFSX1 w2_reg_1__22_ ( .D(n2190), .CK(clk), .SN(rst_n), .Q(n26442), .QN(
        w2[54]) );
  DFFSX1 w2_reg_1__21_ ( .D(n2189), .CK(clk), .SN(rst_n), .Q(n26441), .QN(
        w2[53]) );
  DFFSX1 w2_reg_1__20_ ( .D(n2188), .CK(clk), .SN(rst_n), .Q(n26440), .QN(
        w2[52]) );
  DFFSX1 w2_reg_1__19_ ( .D(n2187), .CK(clk), .SN(rst_n), .Q(n26439), .QN(
        w2[51]) );
  DFFSX1 w2_reg_1__18_ ( .D(n2186), .CK(clk), .SN(rst_n), .Q(n26438), .QN(
        w2[50]) );
  DFFSX1 w2_reg_1__16_ ( .D(n2184), .CK(clk), .SN(rst_n), .Q(n26437), .QN(
        w2[48]) );
  DFFSX1 w2_reg_1__12_ ( .D(n2180), .CK(clk), .SN(rst_n), .Q(n26435), .QN(
        w2[44]) );
  DFFSX1 w2_reg_1__11_ ( .D(n2179), .CK(clk), .SN(rst_n), .Q(n26434), .QN(
        w2[43]) );
  DFFSX1 w2_reg_1__10_ ( .D(n2178), .CK(clk), .SN(rst_n), .Q(n26433), .QN(
        w2[42]) );
  DFFSX1 w2_reg_1__8_ ( .D(n2176), .CK(clk), .SN(rst_n), .Q(n26432), .QN(
        w2[40]) );
  DFFSX1 w2_reg_1__7_ ( .D(n2175), .CK(clk), .SN(rst_n), .Q(n26431), .QN(
        w2[39]) );
  DFFSX1 w2_reg_1__6_ ( .D(n2174), .CK(clk), .SN(rst_n), .Q(n26430), .QN(
        w2[38]) );
  DFFSX1 w2_reg_1__5_ ( .D(n2173), .CK(clk), .SN(rst_n), .Q(n26429), .QN(
        w2[37]) );
  DFFSX1 w2_reg_1__4_ ( .D(n2172), .CK(clk), .SN(rst_n), .Q(n26428), .QN(
        w2[36]) );
  DFFSX1 w2_reg_1__3_ ( .D(n2171), .CK(clk), .SN(rst_n), .Q(n26427), .QN(
        w2[35]) );
  DFFSX1 w2_reg_1__2_ ( .D(n2170), .CK(clk), .SN(rst_n), .Q(n26426), .QN(
        w2[34]) );
  DFFSX1 w2_reg_1__1_ ( .D(n2169), .CK(clk), .SN(rst_n), .Q(n26425), .QN(
        w2[33]) );
  DFFSX1 w2_reg_1__25_ ( .D(n2193), .CK(clk), .SN(rst_n), .Q(n26423), .QN(
        w2[57]) );
  DFFSX1 y20_reg_9_ ( .D(n2369), .CK(clk), .SN(rst_n), .QN(y20[9]) );
  DFFSX1 y20_reg_3_ ( .D(n2363), .CK(clk), .SN(rst_n), .QN(y20[3]) );
  DFFSX1 y20_reg_2_ ( .D(n2362), .CK(clk), .SN(rst_n), .QN(y20[2]) );
  DFFSX1 y20_reg_1_ ( .D(n2361), .CK(clk), .SN(rst_n), .QN(y20[1]) );
  DFFSX1 y20_reg_0_ ( .D(n2360), .CK(clk), .SN(rst_n), .QN(y20[0]) );
  DFFSX1 w2_reg_1__17_ ( .D(n2185), .CK(clk), .SN(rst_n), .Q(n26420), .QN(
        w2[49]) );
  DFFSX1 w2_reg_1__15_ ( .D(n2183), .CK(clk), .SN(rst_n), .Q(n26419), .QN(
        w2[47]) );
  DFFSX1 w2_reg_1__13_ ( .D(n2181), .CK(clk), .SN(rst_n), .Q(n26418), .QN(
        w2[45]) );
  DFFSX1 w2_reg_1__9_ ( .D(n2177), .CK(clk), .SN(rst_n), .Q(n26417), .QN(
        w2[41]) );
  DFFSX1 w2_reg_2__0_ ( .D(n2200), .CK(clk), .SN(rst_n), .QN(w2[64]) );
  DFFSX1 w2_reg_2__29_ ( .D(n2229), .CK(clk), .SN(rst_n), .QN(w2[93]) );
  DFFSX1 w2_reg_2__27_ ( .D(n2227), .CK(clk), .SN(rst_n), .QN(w2[91]) );
  DFFSX1 w2_reg_2__25_ ( .D(n2225), .CK(clk), .SN(rst_n), .QN(w2[89]) );
  DFFSX1 y10_reg_21_ ( .D(n2434), .CK(clk), .SN(rst_n), .Q(n25994), .QN(
        y10[21]) );
  DFFSX1 y10_reg_13_ ( .D(n2418), .CK(clk), .SN(rst_n), .Q(n26222), .QN(
        y10[13]) );
  DFFSX1 y10_reg_7_ ( .D(n2406), .CK(clk), .SN(rst_n), .Q(n26219), .QN(y10[7])
         );
  DFFSX1 y10_reg_3_ ( .D(n2398), .CK(clk), .SN(rst_n), .Q(n25894), .QN(y10[3])
         );
  DFFSX1 y10_reg_16_ ( .D(n2424), .CK(clk), .SN(rst_n), .Q(n26225), .QN(
        y10[16]) );
  DFFSX1 y10_reg_4_ ( .D(n2400), .CK(clk), .SN(rst_n), .Q(n26216), .QN(y10[4])
         );
  DFFSX1 y10_reg_9_ ( .D(n2410), .CK(clk), .SN(rst_n), .Q(n25991), .QN(y10[9])
         );
  DFFSX1 y10_reg_10_ ( .D(n2412), .CK(clk), .SN(rst_n), .Q(n26214), .QN(
        y10[10]) );
  DFFSX1 y10_reg_11_ ( .D(n2414), .CK(clk), .SN(rst_n), .Q(n26215), .QN(
        y10[11]) );
  DFFSX1 y10_reg_29_ ( .D(n2450), .CK(clk), .SN(rst_n), .Q(n26305), .QN(
        y10[29]) );
  DFFSX1 y10_reg_23_ ( .D(n2438), .CK(clk), .SN(rst_n), .Q(n26290), .QN(
        y10[23]) );
  DFFSX1 y10_reg_30_ ( .D(n2452), .CK(clk), .SN(rst_n), .QN(y10[30]) );
  DFFSX1 y10_reg_26_ ( .D(n2444), .CK(clk), .SN(rst_n), .QN(y10[26]) );
  NOR2XL M2_U4_U1_UORT0_1_6 ( .A(M2_b_19_), .B(M2_b_18_), .Y(
        M2_U4_U1_enc_tree_1__1__12_) );
  NAND2XL M2_U3_U1_UOR21_1_2_2 ( .A(M2_U3_U1_enc_tree_1__1__16_), .B(
        M2_U3_U1_enc_tree_1__1__20_), .Y(M2_U3_U1_or2_tree_1__2__16_) );
  NAND2XL M2_U3_U1_UOR21_1_2_3 ( .A(M2_U3_U1_enc_tree_1__1__24_), .B(
        M2_U3_U1_enc_tree_1__1__28_), .Y(M2_U3_U1_or2_tree_1__2__24_) );
  NAND2XL M2_U4_U1_UOR21_1_2_2 ( .A(M2_U4_U1_enc_tree_1__1__16_), .B(
        M2_U4_U1_enc_tree_1__1__20_), .Y(M2_U4_U1_or2_tree_1__2__16_) );
  NAND2XL M2_U4_U1_UOR21_1_2_3 ( .A(M2_U4_U1_enc_tree_1__1__24_), .B(
        M2_U4_U1_enc_tree_1__1__28_), .Y(M2_U4_U1_or2_tree_1__2__24_) );
  NAND2XL M2_U3_U1_UOR21_0_2_2 ( .A(M2_U3_U1_or2_tree_0__1__16_), .B(
        M2_U3_U1_or2_tree_0__1__20_), .Y(M2_U3_U1_or2_tree_0__2__16_) );
  NAND2XL M2_U3_U1_UOR21_0_2_3 ( .A(M2_U3_U1_or2_tree_0__1__24_), .B(
        M2_U3_U1_or2_tree_0__1__28_), .Y(M2_U3_U1_or2_tree_0__2__24_) );
  NAND2XL M2_U4_U1_UOR21_0_2_2 ( .A(M2_U4_U1_or2_tree_0__1__16_), .B(
        M2_U4_U1_or2_tree_0__1__20_), .Y(M2_U4_U1_or2_tree_0__2__16_) );
  NAND2XL M3_U4_U1_UOR21_0_2_2 ( .A(M4_U4_U1_or2_tree_0__1__16_), .B(
        M4_U4_U1_or2_tree_0__1__20_), .Y(M3_U4_U1_or2_tree_0__2__16_) );
  NAND2XL M4_U3_U1_UOR21_0_2_2 ( .A(M4_U3_U1_or2_tree_0__1__16_), .B(
        M4_U3_U1_or2_tree_0__1__20_), .Y(M4_U3_U1_or2_tree_0__2__16_) );
  NAND2XL M4_U3_U1_UOR21_0_2_3 ( .A(M4_U3_U1_or2_tree_0__1__24_), .B(
        M4_U3_U1_or2_tree_0__1__28_), .Y(M4_U3_U1_or2_tree_0__2__24_) );
  NAND2XL M4_U3_U1_UOR21_1_2_2 ( .A(M4_U3_U1_enc_tree_1__1__16_), .B(
        M4_U3_U1_enc_tree_1__1__20_), .Y(M4_U3_U1_or2_tree_1__2__16_) );
  NAND2XL M4_U3_U1_UOR21_1_2_3 ( .A(M4_U3_U1_enc_tree_1__1__24_), .B(
        M4_U3_U1_enc_tree_1__1__28_), .Y(M4_U3_U1_or2_tree_1__2__24_) );
  NAND2XL M3_U3_U1_UOR21_0_2_2 ( .A(M3_U3_U1_or2_tree_0__1__16_), .B(
        M3_U3_U1_or2_tree_0__1__20_), .Y(M3_U3_U1_or2_tree_0__2__16_) );
  NAND2XL M3_U3_U1_UOR21_1_2_2 ( .A(M3_U3_U1_enc_tree_1__1__16_), .B(
        M3_U3_U1_enc_tree_1__1__20_), .Y(M3_U3_U1_or2_tree_1__2__16_) );
  NOR2XL M0_U4_U1_UORT0_1_13 ( .A(M0_b_5_), .B(M0_b_4_), .Y(
        M0_U4_U1_enc_tree_1__1__26_) );
  NOR2XL M0_U4_U1_UORT0_1_11 ( .A(M0_b_9_), .B(M0_b_8_), .Y(
        M0_U4_U1_enc_tree_1__1__22_) );
  NOR2XL M0_U4_U1_UORT0_1_15 ( .A(M0_b_1_), .B(M0_b_0_), .Y(
        M0_U4_U1_enc_tree_1__1__30_) );
  NOR2XL M0_U3_U1_UORT0_1_7 ( .A(n6299), .B(M0_a_16_), .Y(
        M0_U3_U1_enc_tree_1__1__14_) );
  NOR2XL M0_U3_U1_UORT0_1_15 ( .A(n6928), .B(M0_a_0_), .Y(
        M0_U3_U1_enc_tree_1__1__30_) );
  NAND2XL M0_U4_U1_UOR21_0_2_2 ( .A(M0_U4_U1_or2_tree_0__1__16_), .B(
        M0_U4_U1_or2_tree_0__1__20_), .Y(M0_U4_U1_or2_tree_0__2__16_) );
  NAND2XL M0_U3_U1_UOR21_0_2_2 ( .A(M0_U3_U1_or2_tree_0__1__16_), .B(
        M0_U3_U1_or2_tree_0__1__20_), .Y(M0_U3_U1_or2_tree_0__2__16_) );
  NOR2XL M0_U4_U1_UORT0_1_5 ( .A(M0_b_21_), .B(M0_b_20_), .Y(
        M0_U4_U1_enc_tree_1__1__10_) );
  NAND2XL M0_U4_U1_UOR21_1_2_2 ( .A(M0_U4_U1_enc_tree_1__1__16_), .B(
        M0_U4_U1_enc_tree_1__1__20_), .Y(M0_U4_U1_or2_tree_1__2__16_) );
  NOR2XL M0_U3_U1_UORT0_1_5 ( .A(n23219), .B(M0_a_20_), .Y(
        M0_U3_U1_enc_tree_1__1__10_) );
  NAND2XL M0_U3_U1_UOR21_1_2_2 ( .A(M0_U3_U1_enc_tree_1__1__16_), .B(
        M0_U3_U1_enc_tree_1__1__20_), .Y(M0_U3_U1_or2_tree_1__2__16_) );
  NAND2XL M5_U3_U1_UOR21_0_2_2 ( .A(M5_U3_U1_or2_tree_0__1__16_), .B(
        M5_U3_U1_or2_tree_0__1__20_), .Y(M5_U3_U1_or2_tree_0__2__16_) );
  NAND2XL M5_U3_U1_UOR21_1_2_2 ( .A(M5_U3_U1_enc_tree_1__1__16_), .B(
        M5_U3_U1_enc_tree_1__1__20_), .Y(M5_U3_U1_or2_tree_1__2__16_) );
  NOR2XL M1_U4_U1_UORT0_1_15 ( .A(n23174), .B(M1_b_0_), .Y(
        M1_U4_U1_enc_tree_1__1__30_) );
  NOR2XL M1_U3_U1_UORT0_1_12 ( .A(M1_a_7_), .B(M1_a_6_), .Y(
        M1_U3_U1_enc_tree_1__1__24_) );
  NOR2XL M1_U3_U1_UORT0_1_15 ( .A(M1_a_1_), .B(M1_a_0_), .Y(
        M1_U3_U1_enc_tree_1__1__30_) );
  NOR2XL M1_U3_U1_UORT0_1_5 ( .A(M1_a_21_), .B(M1_a_20_), .Y(
        M1_U3_U1_enc_tree_1__1__10_) );
  NAND2XL M1_U3_U1_UOR21_1_2_2 ( .A(M1_U3_U1_enc_tree_1__1__16_), .B(
        M1_U3_U1_enc_tree_1__1__20_), .Y(M1_U3_U1_or2_tree_1__2__16_) );
  NAND2XL M1_U3_U1_UOR21_1_2_3 ( .A(M1_U3_U1_enc_tree_1__1__24_), .B(
        M1_U3_U1_enc_tree_1__1__28_), .Y(M1_U3_U1_or2_tree_1__2__24_) );
  NAND2XL M1_U4_U1_UOR21_1_2_2 ( .A(M1_U4_U1_enc_tree_1__1__16_), .B(
        M1_U4_U1_enc_tree_1__1__20_), .Y(M1_U4_U1_or2_tree_1__2__16_) );
  NAND2XL M1_U4_U1_UOR21_1_2_3 ( .A(M1_U4_U1_enc_tree_1__1__24_), .B(
        M1_U4_U1_enc_tree_1__1__28_), .Y(M1_U4_U1_or2_tree_1__2__24_) );
  NOR2XL M1_U3_U1_UOR20_0_1_4 ( .A(M1_a_15_), .B(M1_a_13_), .Y(
        M1_U3_U1_or2_tree_0__1__16_) );
  NAND2XL M1_U3_U1_UOR21_0_2_2 ( .A(M1_U3_U1_or2_tree_0__1__16_), .B(
        M1_U3_U1_or2_tree_0__1__20_), .Y(M1_U3_U1_or2_tree_0__2__16_) );
  NOR2XL M1_U3_U1_UOR20_0_1_6 ( .A(M1_a_7_), .B(M1_a_5_), .Y(
        M1_U3_U1_or2_tree_0__1__24_) );
  NOR2XL M1_U3_U1_UOR20_0_1_7 ( .A(M1_a_3_), .B(M1_a_1_), .Y(
        M1_U3_U1_or2_tree_0__1__28_) );
  NAND2XL M1_U3_U1_UOR21_0_2_3 ( .A(M1_U3_U1_or2_tree_0__1__24_), .B(
        M1_U3_U1_or2_tree_0__1__28_), .Y(M1_U3_U1_or2_tree_0__2__24_) );
  NAND2XL M1_U4_U1_UOR21_0_2_2 ( .A(M1_U4_U1_or2_tree_0__1__16_), .B(
        M1_U4_U1_or2_tree_0__1__20_), .Y(M1_U4_U1_or2_tree_0__2__16_) );
  NAND2XL M1_U4_U1_UOR21_0_2_3 ( .A(M1_U4_U1_or2_tree_0__1__24_), .B(
        M1_U4_U1_or2_tree_0__1__28_), .Y(M1_U4_U1_or2_tree_0__2__24_) );
  AOI21XL M2_U3_U1_UEN0_0_1_3 ( .A0(M2_a_18_), .A1(n5202), .B0(M2_a_16_), .Y(
        M2_U3_U1_enc_tree_0__1__14_) );
  AOI21XL M2_U3_U1_UEN0_0_1_4 ( .A0(M2_a_14_), .A1(n10338), .B0(M2_a_12_), .Y(
        M2_U3_U1_enc_tree_0__1__18_) );
  AOI21XL M2_U3_U1_UEN0_0_1_6 ( .A0(M2_a_6_), .A1(n9878), .B0(M2_a_4_), .Y(
        M2_U3_U1_enc_tree_0__1__26_) );
  AOI21XL M2_U3_U1_UEN0_0_1_7 ( .A0(M2_a_2_), .A1(n9222), .B0(M2_a_0_), .Y(
        M2_U3_U1_enc_tree_0__1__30_) );
  AOI21XL M2_U4_U1_UEN0_0_1_3 ( .A0(M2_b_18_), .A1(M2_U4_U1_or2_inv_0__14_), 
        .B0(M2_b_16_), .Y(M2_U4_U1_enc_tree_0__1__14_) );
  AOI21XL M2_U4_U1_UEN0_0_1_5 ( .A0(n10342), .A1(M2_U4_U1_or2_inv_0__22_), 
        .B0(M2_b_8_), .Y(M2_U4_U1_enc_tree_0__1__22_) );
  AOI21XL M2_U4_U1_UEN0_0_1_6 ( .A0(M2_b_6_), .A1(M2_U4_U1_or2_inv_0__26_), 
        .B0(M2_b_4_), .Y(M2_U4_U1_enc_tree_0__1__26_) );
  AOI21XL M4_U3_U1_UEN0_0_1_6 ( .A0(M4_a_6_), .A1(n18142), .B0(M4_a_4_), .Y(
        M4_U3_U1_enc_tree_0__1__26_) );
  AOI21XL M3_U3_U1_UEN0_0_1_7 ( .A0(M3_a_2_), .A1(n11691), .B0(n4776), .Y(
        M3_U3_U1_enc_tree_0__1__30_) );
  AOI21XL M0_U3_U1_UEN0_0_1_2 ( .A0(M0_a_22_), .A1(n7711), .B0(M0_a_20_), .Y(
        M0_U3_U1_enc_tree_0__1__10_) );
  AOI21XL M0_U3_U1_UEN0_0_1_3 ( .A0(M0_a_18_), .A1(n7615), .B0(M0_a_16_), .Y(
        M0_U3_U1_enc_tree_0__1__14_) );
  AOI21XL M0_U3_U1_UEN0_0_1_5 ( .A0(M0_a_10_), .A1(n3213), .B0(M0_a_8_), .Y(
        M0_U3_U1_enc_tree_0__1__22_) );
  AOI21XL M0_U3_U1_UEN0_0_1_6 ( .A0(M0_a_6_), .A1(n26488), .B0(M0_a_4_), .Y(
        M0_U3_U1_enc_tree_0__1__26_) );
  AOI21XL M0_U3_U1_UEN0_0_1_7 ( .A0(M0_a_2_), .A1(n6861), .B0(n25871), .Y(
        M0_U3_U1_enc_tree_0__1__30_) );
  AOI21XL M5_U3_U1_UEN0_0_1_2 ( .A0(M5_a_22_), .A1(n6014), .B0(M5_a_20_), .Y(
        M5_U3_U1_enc_tree_0__1__10_) );
  AOI21XL M5_U3_U1_UEN0_0_1_7 ( .A0(M5_a_2_), .A1(n3205), .B0(M5_a_0_), .Y(
        M5_U3_U1_enc_tree_0__1__30_) );
  AOI21XL M1_U3_U1_UEN0_0_1_5 ( .A0(M1_a_10_), .A1(M1_U3_U1_or2_inv_0__22_), 
        .B0(n4565), .Y(M1_U3_U1_enc_tree_0__1__22_) );
  AOI21XL M1_U4_U1_UEN0_0_1_4 ( .A0(M1_b_14_), .A1(n14119), .B0(M1_b_12_), .Y(
        M1_U4_U1_enc_tree_0__1__18_) );
  AOI21XL M1_U4_U1_UEN0_0_1_6 ( .A0(M1_b_6_), .A1(n13842), .B0(M1_b_4_), .Y(
        M1_U4_U1_enc_tree_0__1__26_) );
  AOI21XL M4_U4_U1_UEN0_0_1_2 ( .A0(M3_mult_x_15_b_22_), .A1(
        M4_U4_U1_or2_inv_0__10_), .B0(M3_mult_x_15_b_20_), .Y(
        M4_U4_U1_enc_tree_0__1__10_) );
  DFFSX1 data_reg_2__22_ ( .D(n1700), .CK(clk), .SN(rst_n), .Q(n26265), .QN(
        data[86]) );
  DFFSX1 data_reg_2__13_ ( .D(n1691), .CK(clk), .SN(rst_n), .Q(n26252), .QN(
        data[77]) );
  DFFSX1 data_reg_2__5_ ( .D(n1683), .CK(clk), .SN(rst_n), .QN(data[69]) );
  DFFSX1 data_reg_2__4_ ( .D(n1682), .CK(clk), .SN(rst_n), .QN(data[68]) );
  DFFSX1 data_reg_2__3_ ( .D(n1681), .CK(clk), .SN(rst_n), .Q(n26250), .QN(
        data[67]) );
  DFFSX1 data_reg_2__2_ ( .D(n1680), .CK(clk), .SN(rst_n), .Q(n26267), .QN(
        data[66]) );
  DFFSX1 data_reg_2__1_ ( .D(n1679), .CK(clk), .SN(rst_n), .Q(n26249), .QN(
        data[65]) );
  DFFSX1 data_reg_2__0_ ( .D(n1678), .CK(clk), .SN(rst_n), .Q(n26266), .QN(
        data[64]) );
  DFFSX1 data_reg_1__19_ ( .D(n1665), .CK(clk), .SN(rst_n), .QN(data[51]) );
  DFFSX1 data_reg_1__13_ ( .D(n1659), .CK(clk), .SN(rst_n), .Q(n26259), .QN(
        data[45]) );
  DFFSX1 data_reg_1__4_ ( .D(n1650), .CK(clk), .SN(rst_n), .QN(data[36]) );
  DFFSX1 data_reg_1__2_ ( .D(n1648), .CK(clk), .SN(rst_n), .QN(data[34]) );
  DFFSX1 data_reg_1__1_ ( .D(n1647), .CK(clk), .SN(rst_n), .QN(data[33]) );
  DFFSX1 data_reg_1__0_ ( .D(n1646), .CK(clk), .SN(rst_n), .Q(n26258), .QN(
        data[32]) );
  DFFSX1 data_reg_3__19_ ( .D(n3555), .CK(clk), .SN(rst_n), .Q(n26247), .QN(
        data[115]) );
  DFFSX1 data_reg_3__16_ ( .D(n1726), .CK(clk), .SN(rst_n), .Q(n26024), .QN(
        data[112]) );
  DFFSX1 data_reg_3__15_ ( .D(n1725), .CK(clk), .SN(rst_n), .Q(n26245), .QN(
        data[111]) );
  DFFSX1 data_reg_3__14_ ( .D(n1724), .CK(clk), .SN(rst_n), .Q(n26030), .QN(
        data[110]) );
  DFFSX1 data_reg_3__12_ ( .D(n1722), .CK(clk), .SN(rst_n), .Q(n26279), .QN(
        data[108]) );
  DFFSX1 data_reg_3__7_ ( .D(n1717), .CK(clk), .SN(rst_n), .QN(data[103]) );
  DFFSX1 data_reg_3__22_ ( .D(n1732), .CK(clk), .SN(rst_n), .QN(data[118]) );
  DFFSX1 data_reg_3__2_ ( .D(n1712), .CK(clk), .SN(rst_n), .QN(data[98]) );
  DFFSX1 data_reg_3__17_ ( .D(n1727), .CK(clk), .SN(rst_n), .Q(n26246), .QN(
        data[113]) );
  DFFSX1 data_reg_3__13_ ( .D(n1723), .CK(clk), .SN(rst_n), .Q(n25927), .QN(
        data[109]) );
  DFFSX1 data_reg_3__8_ ( .D(n1718), .CK(clk), .SN(rst_n), .QN(data[104]) );
  DFFSX1 data_reg_3__6_ ( .D(n1716), .CK(clk), .SN(rst_n), .QN(data[102]) );
  DFFSX1 data_reg_3__4_ ( .D(n1714), .CK(clk), .SN(rst_n), .Q(n25933), .QN(
        data[100]) );
  DFFSX1 data_reg_3__3_ ( .D(n1713), .CK(clk), .SN(rst_n), .Q(n26021), .QN(
        data[99]) );
  DFFSX1 data_reg_3__21_ ( .D(n1731), .CK(clk), .SN(rst_n), .QN(data[117]) );
  DFFSX1 data_reg_3__1_ ( .D(n1711), .CK(clk), .SN(rst_n), .QN(data[97]) );
  DFFSX1 data_reg_3__9_ ( .D(n1719), .CK(clk), .SN(rst_n), .QN(data[105]) );
  DFFSX1 data_reg_3__5_ ( .D(n1715), .CK(clk), .SN(rst_n), .Q(n25926), .QN(
        data[101]) );
  DFFSX1 data_reg_3__10_ ( .D(n1720), .CK(clk), .SN(rst_n), .QN(data[106]) );
  DFFSX1 data_reg_3__18_ ( .D(n1728), .CK(clk), .SN(rst_n), .Q(n25928), .QN(
        data[114]) );
  DFFSX1 data_reg_3__11_ ( .D(n1721), .CK(clk), .SN(rst_n), .Q(n26244), .QN(
        data[107]) );
  DFFSX1 data_reg_3__20_ ( .D(n1730), .CK(clk), .SN(rst_n), .Q(n26280), .QN(
        data[116]) );
  DFFSX1 data_reg_3__0_ ( .D(n1710), .CK(clk), .SN(rst_n), .Q(n26288), .QN(
        data[96]) );
  DFFSX1 data_reg_2__21_ ( .D(n1699), .CK(clk), .SN(rst_n), .Q(n2989), .QN(
        data[85]) );
  DFFSX1 data_reg_2__20_ ( .D(n1698), .CK(clk), .SN(rst_n), .Q(n26269), .QN(
        data[84]) );
  DFFSX1 data_reg_2__18_ ( .D(n1696), .CK(clk), .SN(rst_n), .QN(data[82]) );
  DFFSX1 data_reg_2__17_ ( .D(n1695), .CK(clk), .SN(rst_n), .QN(data[81]) );
  DFFSX1 data_reg_2__16_ ( .D(n1694), .CK(clk), .SN(rst_n), .QN(data[80]) );
  DFFSX1 data_reg_2__15_ ( .D(n1693), .CK(clk), .SN(rst_n), .Q(n26253), .QN(
        data[79]) );
  DFFSX1 data_reg_2__14_ ( .D(n1692), .CK(clk), .SN(rst_n), .QN(data[78]) );
  DFFSX1 data_reg_2__11_ ( .D(n1689), .CK(clk), .SN(rst_n), .Q(n26251), .QN(
        data[75]) );
  DFFSX1 data_reg_2__10_ ( .D(n1688), .CK(clk), .SN(rst_n), .QN(data[74]) );
  DFFSX1 data_reg_2__9_ ( .D(n1687), .CK(clk), .SN(rst_n), .QN(data[73]) );
  DFFSX1 data_reg_2__8_ ( .D(n1686), .CK(clk), .SN(rst_n), .QN(data[72]) );
  DFFSX1 data_reg_2__7_ ( .D(n1685), .CK(clk), .SN(rst_n), .QN(data[71]) );
  DFFSX1 data_reg_2__6_ ( .D(n1684), .CK(clk), .SN(rst_n), .QN(data[70]) );
  DFFSX1 data_reg_1__22_ ( .D(n1668), .CK(clk), .SN(rst_n), .Q(n26264), .QN(
        data[54]) );
  DFFSX1 data_reg_1__21_ ( .D(n1667), .CK(clk), .SN(rst_n), .QN(data[53]) );
  DFFSX1 data_reg_1__20_ ( .D(n1666), .CK(clk), .SN(rst_n), .QN(data[52]) );
  DFFSX1 data_reg_1__17_ ( .D(n1663), .CK(clk), .SN(rst_n), .QN(data[49]) );
  DFFSX1 data_reg_1__12_ ( .D(n1658), .CK(clk), .SN(rst_n), .Q(n26242), .QN(
        data[44]) );
  DFFSX1 data_reg_1__11_ ( .D(n1657), .CK(clk), .SN(rst_n), .QN(data[43]) );
  DFFSX1 data_reg_1__10_ ( .D(n1656), .CK(clk), .SN(rst_n), .QN(data[42]) );
  DFFSX1 data_reg_1__9_ ( .D(n1655), .CK(clk), .SN(rst_n), .Q(n26248), .QN(
        data[41]) );
  DFFSX1 data_reg_1__8_ ( .D(n1654), .CK(clk), .SN(rst_n), .Q(n26240), .QN(
        data[40]) );
  DFFSX1 data_reg_1__7_ ( .D(n1653), .CK(clk), .SN(rst_n), .QN(data[39]) );
  DFFSX1 data_reg_1__6_ ( .D(n1652), .CK(clk), .SN(rst_n), .Q(n26239), .QN(
        data[38]) );
  DFFSX1 data_reg_1__5_ ( .D(n1651), .CK(clk), .SN(rst_n), .QN(data[37]) );
  DFFSX1 data_reg_1__3_ ( .D(n1649), .CK(clk), .SN(rst_n), .Q(n26257), .QN(
        data[35]) );
  DFFSX1 iter_reg_5_ ( .D(n1746), .CK(clk), .SN(rst_n), .Q(n26312), .QN(
        iter[5]) );
  DFFSX1 iter_reg_1_ ( .D(n1742), .CK(clk), .SN(rst_n), .Q(n26311), .QN(
        iter[1]) );
  DFFSX1 data_reg_2__19_ ( .D(n1697), .CK(clk), .SN(rst_n), .Q(n26254), .QN(
        data[83]) );
  DFFSX1 data_reg_2__12_ ( .D(n1690), .CK(clk), .SN(rst_n), .QN(data[76]) );
  DFFSX1 data_reg_1__18_ ( .D(n1664), .CK(clk), .SN(rst_n), .Q(n26262), .QN(
        data[50]) );
  DFFSX1 data_reg_1__16_ ( .D(n1662), .CK(clk), .SN(rst_n), .QN(data[48]) );
  DFFSX1 data_reg_1__15_ ( .D(n1661), .CK(clk), .SN(rst_n), .Q(n26261), .QN(
        data[47]) );
  DFFSX1 data_reg_1__14_ ( .D(n1660), .CK(clk), .SN(rst_n), .Q(n26243), .QN(
        data[46]) );
  DFFSX1 w1_reg_3__26_ ( .D(n1858), .CK(clk), .SN(rst_n), .Q(n26328), .QN(
        w1[122]) );
  DFFSX1 w1_reg_3__23_ ( .D(n1846), .CK(clk), .SN(rst_n), .Q(n26329), .QN(
        w1[119]) );
  DFFSX1 w1_reg_3__30_ ( .D(n1874), .CK(clk), .SN(rst_n), .Q(n26351), .QN(
        w1[126]) );
  DFFSX1 w1_reg_3__28_ ( .D(n1866), .CK(clk), .SN(rst_n), .Q(n26331), .QN(
        w1[124]) );
  DFFSX1 w1_reg_3__25_ ( .D(n1854), .CK(clk), .SN(rst_n), .Q(n26330), .QN(
        w1[121]) );
  DFFSX1 w1_reg_2__22_ ( .D(n1841), .CK(clk), .SN(rst_n), .Q(n26093), .QN(
        w1[86]) );
  DFFSX1 w1_reg_1__0_ ( .D(n1752), .CK(clk), .SN(rst_n), .Q(n26354), .QN(
        w1[32]) );
  DFFSX1 w1_reg_6__22_ ( .D(n1969), .CK(clk), .SN(rst_n), .Q(n26076), .QN(
        w1[214]) );
  DFFSX1 w1_reg_6__21_ ( .D(n1965), .CK(clk), .SN(rst_n), .Q(n26082), .QN(
        w1[213]) );
  DFFSX1 w1_reg_4__10_ ( .D(n1923), .CK(clk), .SN(rst_n), .Q(n26062), .QN(
        w1[138]) );
  DFFSX1 w1_reg_3__16_ ( .D(n1818), .CK(clk), .SN(rst_n), .Q(n26339), .QN(
        w1[112]) );
  DFFSX1 w1_reg_3__15_ ( .D(n1814), .CK(clk), .SN(rst_n), .Q(n26340), .QN(
        w1[111]) );
  DFFSX1 w1_reg_3__27_ ( .D(n1862), .CK(clk), .SN(rst_n), .Q(n26332), .QN(
        w1[123]) );
  DFFSX1 w1_reg_2__1_ ( .D(n1757), .CK(clk), .SN(rst_n), .Q(n26098), .QN(
        w1[65]) );
  DFFSX1 w1_reg_6__12_ ( .D(n1929), .CK(clk), .SN(rst_n), .Q(n26074), .QN(
        w1[204]) );
  DFFSX1 w1_reg_4__16_ ( .D(n1947), .CK(clk), .SN(rst_n), .Q(n26066), .QN(
        w1[144]) );
  DFFSX1 w1_reg_5__18_ ( .D(n1952), .CK(clk), .SN(rst_n), .Q(n26319), .QN(
        w1[178]) );
  DFFSX1 w1_reg_6__23_ ( .D(n1973), .CK(clk), .SN(rst_n), .Q(n26099), .QN(
        w1[215]) );
  DFFSX1 w1_reg_5__26_ ( .D(n1984), .CK(clk), .SN(rst_n), .Q(n26322), .QN(
        w1[186]) );
  DFFSX1 w1_reg_1__27_ ( .D(n1860), .CK(clk), .SN(rst_n), .Q(n26352), .QN(
        w1[59]) );
  DFFSX1 w1_reg_1__19_ ( .D(n1828), .CK(clk), .SN(rst_n), .Q(n26326), .QN(
        w1[51]) );
  DFFSX1 w1_reg_4__19_ ( .D(n1959), .CK(clk), .SN(rst_n), .Q(n26065), .QN(
        w1[147]) );
  DFFSX1 w1_reg_6__20_ ( .D(n1961), .CK(clk), .SN(rst_n), .Q(n26083), .QN(
        w1[212]) );
  DFFSX1 w1_reg_6__19_ ( .D(n1957), .CK(clk), .SN(rst_n), .Q(n26077), .QN(
        w1[211]) );
  DFFSX1 w1_reg_2__19_ ( .D(n1829), .CK(clk), .SN(rst_n), .Q(n26054), .QN(
        w1[83]) );
  DFFSX1 w1_reg_1__16_ ( .D(n1816), .CK(clk), .SN(rst_n), .Q(n26104), .QN(
        w1[48]) );
  DFFSX1 w1_reg_6__18_ ( .D(n1953), .CK(clk), .SN(rst_n), .Q(n26050), .QN(
        w1[210]) );
  DFFSX1 w1_reg_6__17_ ( .D(n1949), .CK(clk), .SN(rst_n), .Q(n26084), .QN(
        w1[209]) );
  DFFSX1 w1_reg_2__18_ ( .D(n1825), .CK(clk), .SN(rst_n), .Q(n26094), .QN(
        w1[82]) );
  DFFSX1 w1_reg_5__30_ ( .D(n2000), .CK(clk), .SN(rst_n), .Q(n26325), .QN(
        w1[190]) );
  DFFSX1 w1_reg_0__17_ ( .D(n1823), .CK(clk), .SN(rst_n), .Q(n26071), .QN(
        w1[17]) );
  DFFSX1 w1_reg_7__10_ ( .D(n1922), .CK(clk), .SN(rst_n), .Q(n26390), .QN(
        w1[234]) );
  DFFSX1 w1_reg_7__8_ ( .D(n1914), .CK(clk), .SN(rst_n), .Q(n26392), .QN(
        w1[232]) );
  DFFSX1 w1_reg_7__12_ ( .D(n1930), .CK(clk), .SN(rst_n), .Q(n26388), .QN(
        w1[236]) );
  DFFSX1 w1_reg_7__11_ ( .D(n1926), .CK(clk), .SN(rst_n), .Q(n26389), .QN(
        w1[235]) );
  DFFSX1 w1_reg_7__7_ ( .D(n1910), .CK(clk), .SN(rst_n), .Q(n26393), .QN(
        w1[231]) );
  DFFSX1 w1_reg_7__5_ ( .D(n1902), .CK(clk), .SN(rst_n), .Q(n26395), .QN(
        w1[229]) );
  DFFSX1 w1_reg_7__18_ ( .D(n1954), .CK(clk), .SN(rst_n), .Q(n26383), .QN(
        w1[242]) );
  DFFSX1 w1_reg_7__17_ ( .D(n1950), .CK(clk), .SN(rst_n), .Q(n26384), .QN(
        w1[241]) );
  DFFSX1 w1_reg_7__15_ ( .D(n1942), .CK(clk), .SN(rst_n), .Q(n26385), .QN(
        w1[239]) );
  DFFSX1 w1_reg_7__14_ ( .D(n1938), .CK(clk), .SN(rst_n), .Q(n26386), .QN(
        w1[238]) );
  DFFSX1 w1_reg_7__13_ ( .D(n1934), .CK(clk), .SN(rst_n), .Q(n26387), .QN(
        w1[237]) );
  DFFSX1 w1_reg_3__18_ ( .D(n1826), .CK(clk), .SN(rst_n), .Q(n26404), .QN(
        w1[114]) );
  DFFSX1 w1_reg_7__2_ ( .D(n1890), .CK(clk), .SN(rst_n), .Q(n26398), .QN(
        w1[226]) );
  DFFSX1 w1_reg_7__1_ ( .D(n1886), .CK(clk), .SN(rst_n), .Q(n26399), .QN(
        w1[225]) );
  DFFSX1 w1_reg_3__1_ ( .D(n1758), .CK(clk), .SN(rst_n), .Q(n26408), .QN(
        w1[97]) );
  DFFSX1 w1_reg_7__30_ ( .D(n2002), .CK(clk), .SN(rst_n), .Q(n26401), .QN(
        w1[254]) );
  DFFSX1 w1_reg_7__26_ ( .D(n1986), .CK(clk), .SN(rst_n), .Q(n26371), .QN(
        w1[250]) );
  DFFSX1 w1_reg_3__0_ ( .D(n1754), .CK(clk), .SN(rst_n), .Q(n26409), .QN(
        w1[96]) );
  DFFSX1 w1_reg_7__4_ ( .D(n1898), .CK(clk), .SN(rst_n), .Q(n26396), .QN(
        w1[228]) );
  DFFSX1 w1_reg_7__0_ ( .D(n1882), .CK(clk), .SN(rst_n), .Q(n26400), .QN(
        w1[224]) );
  DFFSX1 w1_reg_7__9_ ( .D(n1918), .CK(clk), .SN(rst_n), .Q(n26391), .QN(
        w1[233]) );
  DFFSX1 w1_reg_3__5_ ( .D(n1774), .CK(clk), .SN(rst_n), .Q(n26406), .QN(
        w1[101]) );
  DFFSX1 w1_reg_7__6_ ( .D(n1906), .CK(clk), .SN(rst_n), .Q(n26394), .QN(
        w1[230]) );
  DFFSX1 w1_reg_3__6_ ( .D(n1778), .CK(clk), .SN(rst_n), .Q(n26405), .QN(
        w1[102]) );
  DFFSX1 w1_reg_7__3_ ( .D(n1894), .CK(clk), .SN(rst_n), .Q(n26397), .QN(
        w1[227]) );
  DFFSX1 w1_reg_3__4_ ( .D(n1770), .CK(clk), .SN(rst_n), .Q(n26407), .QN(
        w1[100]) );
  DFFSX1 w1_reg_7__21_ ( .D(n1966), .CK(clk), .SN(rst_n), .Q(n26380), .QN(
        w1[245]) );
  DFFSX1 w1_reg_7__20_ ( .D(n1962), .CK(clk), .SN(rst_n), .Q(n26381), .QN(
        w1[244]) );
  DFFSX1 w1_reg_7__22_ ( .D(n1970), .CK(clk), .SN(rst_n), .Q(n26379), .QN(
        w1[246]) );
  DFFSX1 w1_reg_7__31_ ( .D(n2006), .CK(clk), .SN(rst_n), .Q(n26378), .QN(
        w1[255]) );
  DFFSX1 w1_reg_3__22_ ( .D(n1842), .CK(clk), .SN(rst_n), .Q(n26402), .QN(
        w1[118]) );
  DFFSX1 w1_reg_7__24_ ( .D(n1978), .CK(clk), .SN(rst_n), .Q(n26376), .QN(
        w1[248]) );
  DFFSX1 w1_reg_3__19_ ( .D(n1830), .CK(clk), .SN(rst_n), .Q(n26403), .QN(
        w1[115]) );
  DFFSX1 w1_reg_7__19_ ( .D(n1958), .CK(clk), .SN(rst_n), .Q(n26382), .QN(
        w1[243]) );
  DFFSX1 w1_reg_7__23_ ( .D(n1974), .CK(clk), .SN(rst_n), .Q(n26372), .QN(
        w1[247]) );
  DFFSX1 w1_reg_7__29_ ( .D(n1998), .CK(clk), .SN(rst_n), .Q(n26375), .QN(
        w1[253]) );
  DFFSX1 w1_reg_7__27_ ( .D(n1990), .CK(clk), .SN(rst_n), .Q(n26374), .QN(
        w1[251]) );
  DFFSX1 w1_reg_7__25_ ( .D(n1982), .CK(clk), .SN(rst_n), .Q(n26373), .QN(
        w1[249]) );
  DFFSX1 w1_reg_2__5_ ( .D(n1773), .CK(clk), .SN(rst_n), .Q(n26096), .QN(
        w1[69]) );
  DFFSX1 w1_reg_6__29_ ( .D(n1997), .CK(clk), .SN(rst_n), .Q(n26101), .QN(
        w1[221]) );
  DFFSX1 w1_reg_6__27_ ( .D(n1989), .CK(clk), .SN(rst_n), .Q(n26056), .QN(
        w1[219]) );
  DFFSX1 w1_reg_5__27_ ( .D(n1988), .CK(clk), .SN(rst_n), .Q(n26323), .QN(
        w1[187]) );
  DFFSX1 w1_reg_0__27_ ( .D(n1863), .CK(clk), .SN(rst_n), .Q(n26069), .QN(
        w1[27]) );
  DFFSX1 w1_reg_6__5_ ( .D(n1901), .CK(clk), .SN(rst_n), .Q(n26079), .QN(
        w1[197]) );
  DFFSX1 w1_reg_6__28_ ( .D(n1993), .CK(clk), .SN(rst_n), .Q(n26100), .QN(
        w1[220]) );
  DFFSX1 w1_reg_6__26_ ( .D(n1985), .CK(clk), .SN(rst_n), .Q(n26055), .QN(
        w1[218]) );
  DFFSX1 w1_reg_6__25_ ( .D(n1981), .CK(clk), .SN(rst_n), .Q(n26057), .QN(
        w1[217]) );
  DFFSX1 w1_reg_6__9_ ( .D(n1917), .CK(clk), .SN(rst_n), .Q(n26089), .QN(
        w1[201]) );
  DFFSX1 w1_reg_6__8_ ( .D(n1913), .CK(clk), .SN(rst_n), .Q(n26090), .QN(
        w1[200]) );
  DFFSX1 w1_reg_4__9_ ( .D(n1919), .CK(clk), .SN(rst_n), .Q(n26063), .QN(
        w1[137]) );
  DFFSX1 w1_reg_4__8_ ( .D(n1915), .CK(clk), .SN(rst_n), .Q(n26064), .QN(
        w1[136]) );
  DFFSX1 w1_reg_5__0_ ( .D(n1880), .CK(clk), .SN(rst_n), .Q(n26317), .QN(
        w1[160]) );
  DFFSX1 w1_reg_3__24_ ( .D(n1850), .CK(clk), .SN(rst_n), .Q(n26334), .QN(
        w1[120]) );
  DFFSX1 w1_reg_3__21_ ( .D(n1838), .CK(clk), .SN(rst_n), .Q(n26336), .QN(
        w1[117]) );
  DFFSX1 w1_reg_3__17_ ( .D(n1822), .CK(clk), .SN(rst_n), .Q(n26338), .QN(
        w1[113]) );
  DFFSX1 w1_reg_3__10_ ( .D(n1794), .CK(clk), .SN(rst_n), .Q(n26345), .QN(
        w1[106]) );
  DFFSX1 w1_reg_3__9_ ( .D(n1790), .CK(clk), .SN(rst_n), .Q(n26346), .QN(
        w1[105]) );
  DFFSX1 w1_reg_3__7_ ( .D(n1782), .CK(clk), .SN(rst_n), .Q(n26348), .QN(
        w1[103]) );
  DFFSX1 w1_reg_3__31_ ( .D(n1878), .CK(clk), .SN(rst_n), .Q(n26335), .QN(
        w1[127]) );
  DFFSX1 w1_reg_3__14_ ( .D(n1810), .CK(clk), .SN(rst_n), .Q(n26341), .QN(
        w1[110]) );
  DFFSX1 w1_reg_3__13_ ( .D(n1806), .CK(clk), .SN(rst_n), .Q(n26342), .QN(
        w1[109]) );
  DFFSX1 w1_reg_7__16_ ( .D(n1946), .CK(clk), .SN(rst_n), .Q(n26327), .QN(
        w1[240]) );
  DFFSX1 w1_reg_3__29_ ( .D(n1870), .CK(clk), .SN(rst_n), .Q(n26333), .QN(
        w1[125]) );
  DFFSX1 w1_reg_2__10_ ( .D(n1793), .CK(clk), .SN(rst_n), .Q(n26363), .QN(
        w1[74]) );
  DFFSX1 w1_reg_4__31_ ( .D(n2007), .CK(clk), .SN(rst_n), .Q(n26313), .QN(
        w1[159]) );
  DFFSX1 w1_reg_1__5_ ( .D(n1772), .CK(clk), .SN(rst_n), .Q(n26366), .QN(
        w1[37]) );
  DFFSX1 w1_reg_1__3_ ( .D(n1764), .CK(clk), .SN(rst_n), .Q(n26367), .QN(
        w1[35]) );
  DFFSX1 w1_reg_1__2_ ( .D(n1760), .CK(clk), .SN(rst_n), .Q(n26368), .QN(
        w1[34]) );
  DFFSX1 w1_reg_1__29_ ( .D(n1868), .CK(clk), .SN(rst_n), .Q(n26353), .QN(
        w1[61]) );
  DFFSX1 w1_reg_5__10_ ( .D(n1920), .CK(clk), .SN(rst_n), .Q(n26358), .QN(
        w1[170]) );
  DFFSX1 w1_reg_5__9_ ( .D(n1916), .CK(clk), .SN(rst_n), .Q(n26359), .QN(
        w1[169]) );
  DFFSX1 w1_reg_5__8_ ( .D(n1912), .CK(clk), .SN(rst_n), .Q(n26360), .QN(
        w1[168]) );
  DFFSX1 w1_reg_2__12_ ( .D(n1801), .CK(clk), .SN(rst_n), .Q(n26362), .QN(
        w1[76]) );
  DFFSX1 w1_reg_1__14_ ( .D(n1808), .CK(clk), .SN(rst_n), .Q(n26365), .QN(
        w1[46]) );
  DFFSX1 w1_reg_0__9_ ( .D(n1791), .CK(clk), .SN(rst_n), .Q(n26260), .QN(w1[9]) );
  DFFSX1 w1_reg_0__1_ ( .D(n1759), .CK(clk), .SN(rst_n), .Q(n26287), .QN(w1[1]) );
  DFFSX1 w1_reg_3__20_ ( .D(n1834), .CK(clk), .SN(rst_n), .Q(n26337), .QN(
        w1[116]) );
  DFFSX1 w1_reg_3__12_ ( .D(n1802), .CK(clk), .SN(rst_n), .Q(n26343), .QN(
        w1[108]) );
  DFFSX1 w1_reg_3__11_ ( .D(n1798), .CK(clk), .SN(rst_n), .Q(n26344), .QN(
        w1[107]) );
  DFFSX1 w1_reg_3__8_ ( .D(n1786), .CK(clk), .SN(rst_n), .Q(n26347), .QN(
        w1[104]) );
  DFFSX1 w1_reg_3__2_ ( .D(n1762), .CK(clk), .SN(rst_n), .Q(n26350), .QN(
        w1[98]) );
  DFFSX1 w1_reg_3__3_ ( .D(n1766), .CK(clk), .SN(rst_n), .Q(n26349), .QN(
        w1[99]) );
  DFFSX1 w1_reg_2__0_ ( .D(n1753), .CK(clk), .SN(rst_n), .Q(n26075), .QN(
        w1[64]) );
  DFFSX1 w1_reg_6__14_ ( .D(n1937), .CK(clk), .SN(rst_n), .Q(n26086), .QN(
        w1[206]) );
  DFFSX1 w1_reg_6__13_ ( .D(n1933), .CK(clk), .SN(rst_n), .Q(n26051), .QN(
        w1[205]) );
  DFFSX1 w1_reg_6__30_ ( .D(n2001), .CK(clk), .SN(rst_n), .Q(n26059), .QN(
        w1[222]) );
  DFFSX1 w1_reg_0__0_ ( .D(n1755), .CK(clk), .SN(rst_n), .Q(n26068), .QN(w1[0]) );
  DFFSX1 w1_reg_2__6_ ( .D(n1777), .CK(clk), .SN(rst_n), .Q(n26095), .QN(
        w1[70]) );
  DFFSX1 w1_reg_7__28_ ( .D(n1994), .CK(clk), .SN(rst_n), .Q(n26355), .QN(
        w1[252]) );
  DFFSX1 w1_reg_6__3_ ( .D(n1893), .CK(clk), .SN(rst_n), .Q(n26092), .QN(
        w1[195]) );
  DFFSX1 w1_reg_6__2_ ( .D(n1889), .CK(clk), .SN(rst_n), .Q(n26052), .QN(
        w1[194]) );
  DFFSX1 w1_reg_1__10_ ( .D(n1792), .CK(clk), .SN(rst_n), .Q(n26105), .QN(
        w1[42]) );
  DFFSX1 w1_reg_6__31_ ( .D(n2005), .CK(clk), .SN(rst_n), .Q(n26103), .QN(
        w1[223]) );
  DFFSX1 w1_reg_6__15_ ( .D(n1941), .CK(clk), .SN(rst_n), .Q(n26085), .QN(
        w1[207]) );
  DFFSX1 w1_reg_6__11_ ( .D(n1925), .CK(clk), .SN(rst_n), .Q(n26087), .QN(
        w1[203]) );
  DFFSX1 w1_reg_6__10_ ( .D(n1921), .CK(clk), .SN(rst_n), .Q(n26088), .QN(
        w1[202]) );
  DFFSX1 w1_reg_0__14_ ( .D(n1811), .CK(clk), .SN(rst_n), .Q(n26072), .QN(
        w1[14]) );
  DFFSX1 w1_reg_6__24_ ( .D(n1977), .CK(clk), .SN(rst_n), .Q(n26102), .QN(
        w1[216]) );
  DFFSX1 w1_reg_6__7_ ( .D(n1909), .CK(clk), .SN(rst_n), .Q(n26091), .QN(
        w1[199]) );
  DFFSX1 w1_reg_6__6_ ( .D(n1905), .CK(clk), .SN(rst_n), .Q(n26078), .QN(
        w1[198]) );
  DFFSX1 w1_reg_5__25_ ( .D(n1980), .CK(clk), .SN(rst_n), .Q(n26324), .QN(
        w1[185]) );
  DFFSX1 w1_reg_0__29_ ( .D(n1871), .CK(clk), .SN(rst_n), .Q(n26070), .QN(
        w1[29]) );
  DFFSX1 w1_reg_6__4_ ( .D(n1897), .CK(clk), .SN(rst_n), .Q(n26080), .QN(
        w1[196]) );
  DFFSX1 w1_reg_1__12_ ( .D(n1800), .CK(clk), .SN(rst_n), .Q(n26058), .QN(
        w1[44]) );
  DFFSX1 w1_reg_5__13_ ( .D(n1932), .CK(clk), .SN(rst_n), .Q(n26320), .QN(
        w1[173]) );
  DFFSX1 w1_reg_0__12_ ( .D(n1803), .CK(clk), .SN(rst_n), .Q(n26315), .QN(
        w1[12]) );
  DFFSX1 w1_reg_6__1_ ( .D(n1885), .CK(clk), .SN(rst_n), .Q(n26081), .QN(
        w1[193]) );
  DFFSX1 w1_reg_6__0_ ( .D(n1881), .CK(clk), .SN(rst_n), .Q(n26053), .QN(
        w1[192]) );
  DFFSX1 w1_reg_5__2_ ( .D(n1888), .CK(clk), .SN(rst_n), .Q(n26321), .QN(
        w1[162]) );
  DFFSX1 w1_reg_0__2_ ( .D(n1763), .CK(clk), .SN(rst_n), .Q(n26027), .QN(w1[2]) );
  DFFSX1 w1_reg_2__4_ ( .D(n1769), .CK(clk), .SN(rst_n), .Q(n26097), .QN(
        w1[68]) );
  DFFSX1 w1_reg_0__3_ ( .D(n1767), .CK(clk), .SN(rst_n), .Q(n26039), .QN(w1[3]) );
  DFFSX1 w1_reg_0__5_ ( .D(n1775), .CK(clk), .SN(rst_n), .Q(n26073), .QN(w1[5]) );
  DFFSX1 w1_reg_2__16_ ( .D(n1817), .CK(clk), .SN(rst_n), .Q(n26361), .QN(
        w1[80]) );
  DFFSX1 w1_reg_5__16_ ( .D(n1944), .CK(clk), .SN(rst_n), .Q(n26357), .QN(
        w1[176]) );
  DFFSX1 w1_reg_5__19_ ( .D(n1956), .CK(clk), .SN(rst_n), .Q(n26356), .QN(
        w1[179]) );
  DFFSX1 w1_reg_1__17_ ( .D(n1820), .CK(clk), .SN(rst_n), .Q(n26364), .QN(
        w1[49]) );
  DFFSX1 sigma12_reg_31_ ( .D(n2358), .CK(clk), .SN(rst_n), .Q(n26316), .QN(
        sigma12[31]) );
  DFFSX1 sigma11_reg_31_ ( .D(n2359), .CK(clk), .SN(rst_n), .Q(n26067), .QN(
        sigma11[31]) );
  DFFSX1 sigma10_reg_31_ ( .D(n2295), .CK(clk), .SN(rst_n), .Q(n26310), .QN(
        sigma10[31]) );
  DFFSX1 target_temp_reg_31_ ( .D(n2263), .CK(clk), .SN(rst_n), .Q(n25992), 
        .QN(target_temp[31]) );
  DFFSX1 w1_reg_10__31_ ( .D(n2133), .CK(clk), .SN(rst_n), .Q(n26049), .QN(
        w1[351]) );
  DFFSX1 w2_reg_1__31_ ( .D(n2199), .CK(clk), .SN(rst_n), .Q(n26314), .QN(
        w2[63]) );
  DFFSX1 y11_reg_31_ ( .D(n2487), .CK(clk), .SN(rst_n), .Q(n26195), .QN(
        y11[31]) );
  DFFSX1 y12_reg_31_ ( .D(n2455), .CK(clk), .SN(rst_n), .Q(n26227), .QN(
        y12[31]) );
  DFFSX1 w1_reg_11__31_ ( .D(n2134), .CK(clk), .SN(rst_n), .Q(n26377), .QN(
        w1[383]) );
  DFFSX1 w2_reg_0__31_ ( .D(n2167), .CK(clk), .SN(rst_n), .Q(n26048), .QN(
        w2[31]) );
  DFFSX1 w1_reg_9__31_ ( .D(n2132), .CK(clk), .SN(rst_n), .Q(n26318), .QN(
        w1[319]) );
  DFFSX1 y10_reg_31_ ( .D(n2454), .CK(clk), .SN(rst_n), .Q(n26213), .QN(
        y10[31]) );
  DFFSX1 target_temp_reg_9_ ( .D(n2241), .CK(clk), .SN(rst_n), .Q(n25888), 
        .QN(target_temp[9]) );
  DFFSX1 target_temp_reg_2_ ( .D(n2234), .CK(clk), .SN(rst_n), .Q(n26256), 
        .QN(target_temp[2]) );
  DFFSX1 target_temp_reg_3_ ( .D(n2235), .CK(clk), .SN(rst_n), .Q(n26255), 
        .QN(target_temp[3]) );
  DFFSX1 target_temp_reg_1_ ( .D(n2233), .CK(clk), .SN(rst_n), .Q(n26025), 
        .QN(target_temp[1]) );
  DFFSX1 target_temp_reg_22_ ( .D(n2254), .CK(clk), .SN(rst_n), .Q(n26141), 
        .QN(target_temp[22]) );
  DFFSX1 target_temp_reg_29_ ( .D(n2261), .CK(clk), .SN(rst_n), .Q(n26144), 
        .QN(target_temp[29]) );
  DFFSX1 target_temp_reg_26_ ( .D(n2258), .CK(clk), .SN(rst_n), .Q(n26145), 
        .QN(target_temp[26]) );
  DFFSX1 target_temp_reg_25_ ( .D(n2257), .CK(clk), .SN(rst_n), .Q(n26143), 
        .QN(target_temp[25]) );
  DFFSX1 w1_reg_10__30_ ( .D(n2129), .CK(clk), .SN(rst_n), .Q(n26134), .QN(
        w1[350]) );
  DFFSX1 w1_reg_10__29_ ( .D(n2125), .CK(clk), .SN(rst_n), .Q(n26113), .QN(
        w1[349]) );
  DFFSX1 w1_reg_10__28_ ( .D(n2121), .CK(clk), .SN(rst_n), .Q(n26112), .QN(
        w1[348]) );
  DFFSX1 w1_reg_10__24_ ( .D(n2105), .CK(clk), .SN(rst_n), .Q(n26114), .QN(
        w1[344]) );
  DFFSX1 w1_reg_10__23_ ( .D(n2101), .CK(clk), .SN(rst_n), .Q(n26110), .QN(
        w1[343]) );
  DFFSX1 w1_reg_10__26_ ( .D(n2113), .CK(clk), .SN(rst_n), .Q(n26109), .QN(
        w1[346]) );
  DFFSX1 w1_reg_10__25_ ( .D(n2109), .CK(clk), .SN(rst_n), .Q(n26111), .QN(
        w1[345]) );
  DFFSX1 w1_reg_10__4_ ( .D(n2025), .CK(clk), .SN(rst_n), .Q(n26129), .QN(
        w1[324]) );
  DFFSX1 w1_reg_10__5_ ( .D(n2029), .CK(clk), .SN(rst_n), .Q(n26128), .QN(
        w1[325]) );
  DFFSX1 w2_reg_1__27_ ( .D(n2195), .CK(clk), .SN(rst_n), .Q(n26421), .QN(
        w2[59]) );
  DFFSX1 w1_reg_10__7_ ( .D(n2037), .CK(clk), .SN(rst_n), .Q(n26126), .QN(
        w1[327]) );
  DFFSX1 w1_reg_10__16_ ( .D(n2073), .CK(clk), .SN(rst_n), .Q(n26135), .QN(
        w1[336]) );
  DFFSX1 w1_reg_10__6_ ( .D(n2033), .CK(clk), .SN(rst_n), .Q(n26127), .QN(
        w1[326]) );
  DFFSX1 w2_reg_1__30_ ( .D(n2198), .CK(clk), .SN(rst_n), .Q(n26304), .QN(
        w2[62]) );
  DFFSX1 w2_reg_1__29_ ( .D(n2197), .CK(clk), .SN(rst_n), .Q(n26422), .QN(
        w2[61]) );
  DFFSX1 w2_reg_1__28_ ( .D(n2196), .CK(clk), .SN(rst_n), .Q(n26044), .QN(
        w2[60]) );
  DFFXL temp3_reg_24_ ( .D(mul5_out[24]), .CK(clk), .Q(temp3[24]) );
  DFFSX4 y20_reg_22_ ( .D(n2382), .CK(clk), .SN(rst_n), .Q(n26169), .QN(
        y20[22]) );
  DFFXL temp0_reg_28_ ( .D(n2560), .CK(clk), .Q(temp0[28]), .QN(n26514) );
  DFFXL temp0_reg_27_ ( .D(n2562), .CK(clk), .Q(temp0[27]), .QN(n26515) );
  DFFXL temp0_reg_29_ ( .D(n2558), .CK(clk), .Q(temp0[29]), .QN(n26594) );
  DFFXL temp0_reg_26_ ( .D(n2564), .CK(clk), .Q(temp0[26]), .QN(n26546) );
  DFFXL temp0_reg_24_ ( .D(n2568), .CK(clk), .Q(temp0[24]), .QN(n26545) );
  DFFXL temp3_reg_9_ ( .D(mul5_out[9]), .CK(clk), .Q(temp3[9]) );
  DFFXL temp3_reg_8_ ( .D(mul5_out[8]), .CK(clk), .Q(temp3[8]) );
  DFFXL temp3_reg_5_ ( .D(mul5_out[5]), .CK(clk), .Q(temp3[5]) );
  DFFXL temp3_reg_4_ ( .D(mul5_out[4]), .CK(clk), .Q(temp3[4]) );
  DFFXL temp0_reg_21_ ( .D(n2574), .CK(clk), .Q(temp0[21]), .QN(n26572) );
  DFFXL temp0_reg_20_ ( .D(n2576), .CK(clk), .Q(temp0[20]), .QN(n26573) );
  DFFXL temp2_reg_1_ ( .D(n2615), .CK(clk), .Q(temp2[1]), .QN(n26543) );
  DFFXL temp2_reg_16_ ( .D(n2585), .CK(clk), .Q(temp2[16]), .QN(n26526) );
  DFFXL temp3_reg_0_ ( .D(mul5_out[0]), .CK(clk), .Q(temp3[0]) );
  DFFXL temp2_reg_0_ ( .D(n2617), .CK(clk), .Q(temp2[0]), .QN(n26544) );
  DFFXL temp2_reg_19_ ( .D(n2579), .CK(clk), .Q(temp2[19]), .QN(n26523) );
  DFFXL temp0_reg_4_ ( .D(n2608), .CK(clk), .Q(temp0[4]), .QN(n26589) );
  DFFXL temp2_reg_20_ ( .D(n2577), .CK(clk), .Q(temp2[20]), .QN(n26522) );
  DFFXL temp1_reg_23_ ( .D(n2531), .CK(clk), .Q(temp1[23]), .QN(n26509) );
  DFFXL temp1_reg_30_ ( .D(n2524), .CK(clk), .Q(temp1[30]), .QN(n26507) );
  DFFXL temp1_reg_27_ ( .D(n2527), .CK(clk), .Q(temp1[27]), .QN(n26512) );
  DFFXL temp1_reg_26_ ( .D(n2528), .CK(clk), .Q(temp1[26]), .QN(n26505) );
  DFFXL temp1_reg_25_ ( .D(n2529), .CK(clk), .Q(temp1[25]), .QN(n26511) );
  DFFXL temp1_reg_24_ ( .D(n2530), .CK(clk), .Q(temp1[24]), .QN(n26510) );
  DFFXL temp1_reg_29_ ( .D(n2525), .CK(clk), .Q(temp1[29]), .QN(n26508) );
  DFFXL temp1_reg_28_ ( .D(n2526), .CK(clk), .Q(temp1[28]), .QN(n26506) );
  DFFXL temp1_reg_2_ ( .D(n2552), .CK(clk), .Q(temp1[2]), .QN(n26568) );
  DFFXL temp1_reg_15_ ( .D(n2539), .CK(clk), .Q(temp1[15]), .QN(n26555) );
  DFFXL temp3_reg_17_ ( .D(mul5_out[17]), .CK(clk), .Q(temp3[17]) );
  DFFXL temp1_reg_17_ ( .D(n2537), .CK(clk), .Q(temp1[17]), .QN(n26553) );
  DFFXL temp1_reg_19_ ( .D(n2535), .CK(clk), .Q(temp1[19]), .QN(n26551) );
  DFFXL temp2_reg_15_ ( .D(n2587), .CK(clk), .Q(temp2[15]), .QN(n26527) );
  DFFXL temp2_reg_10_ ( .D(n2597), .CK(clk), .Q(temp2[10]), .QN(n26532) );
  DFFXL temp2_reg_8_ ( .D(n2601), .CK(clk), .Q(temp2[8]), .QN(n26535) );
  DFFXL temp2_reg_6_ ( .D(n2605), .CK(clk), .Q(temp2[6]), .QN(n26538) );
  DFFXL temp2_reg_3_ ( .D(n2611), .CK(clk), .Q(temp2[3]), .QN(n26541) );
  DFFXL temp1_reg_20_ ( .D(n2534), .CK(clk), .Q(temp1[20]), .QN(n26550) );
  DFFXL temp2_reg_2_ ( .D(n2613), .CK(clk), .Q(temp2[2]), .QN(n26542) );
  DFFXL temp0_reg_22_ ( .D(n2572), .CK(clk), .Q(temp0[22]), .QN(n26571) );
  DFFXL temp3_reg_2_ ( .D(mul5_out[2]), .CK(clk), .Q(temp3[2]) );
  DFFXL temp1_reg_11_ ( .D(n2543), .CK(clk), .Q(temp1[11]), .QN(n26559) );
  DFFXL temp2_reg_17_ ( .D(n2583), .CK(clk), .Q(temp2[17]), .QN(n26525) );
  DFFXL temp2_reg_30_ ( .D(n2557), .CK(clk), .Q(temp2[30]), .QN(n26497) );
  DFFXL temp1_reg_6_ ( .D(n2548), .CK(clk), .Q(temp1[6]), .QN(n26564) );
  DFFXL temp3_reg_16_ ( .D(mul5_out[16]), .CK(clk), .Q(temp3[16]) );
  DFFXL temp1_reg_0_ ( .D(n2554), .CK(clk), .Q(temp1[0]), .QN(n26570) );
  DFFXL temp3_reg_14_ ( .D(mul5_out[14]), .CK(clk), .Q(temp3[14]) );
  DFFXL temp3_reg_7_ ( .D(mul5_out[7]), .CK(clk), .Q(temp3[7]) );
  DFFXL temp3_reg_3_ ( .D(mul5_out[3]), .CK(clk), .Q(temp3[3]) );
  DFFXL temp1_reg_4_ ( .D(n2550), .CK(clk), .Q(temp1[4]), .QN(n26566) );
  DFFXL temp1_reg_1_ ( .D(n2553), .CK(clk), .Q(temp1[1]), .QN(n26569) );
  DFFXL temp0_reg_1_ ( .D(n2614), .CK(clk), .Q(temp0[1]), .QN(n26592) );
  DFFXL temp3_reg_15_ ( .D(mul5_out[15]), .CK(clk), .Q(temp3[15]) );
  DFFXL temp3_reg_22_ ( .D(mul5_out[22]), .CK(clk), .Q(temp3[22]) );
  DFFXL temp3_reg_6_ ( .D(mul5_out[6]), .CK(clk), .Q(temp3[6]) );
  DFFXL temp1_reg_8_ ( .D(n2546), .CK(clk), .Q(temp1[8]), .QN(n26562) );
  DFFXL temp0_reg_0_ ( .D(n2616), .CK(clk), .Q(temp0[0]), .QN(n26593) );
  DFFXL temp0_reg_13_ ( .D(n2590), .CK(clk), .Q(temp0[13]), .QN(n26580) );
  DFFXL temp3_reg_1_ ( .D(mul5_out[1]), .CK(clk), .Q(temp3[1]) );
  DFFXL temp0_reg_2_ ( .D(n2612), .CK(clk), .Q(temp0[2]), .QN(n26591) );
  DFFXL temp2_reg_23_ ( .D(n2571), .CK(clk), .Q(temp2[23]), .QN(n26500) );
  DFFXL temp3_reg_18_ ( .D(mul5_out[18]), .CK(clk), .Q(temp3[18]) );
  DFFXL temp1_reg_22_ ( .D(n2532), .CK(clk), .Q(temp1[22]), .QN(n26548) );
  DFFXL temp1_reg_7_ ( .D(n2547), .CK(clk), .Q(temp1[7]), .QN(n26563) );
  DFFXL temp2_reg_13_ ( .D(n2591), .CK(clk), .Q(temp2[13]), .QN(n26529) );
  DFFXL temp2_reg_11_ ( .D(n2595), .CK(clk), .Q(temp2[11]), .QN(n26531) );
  DFFXL temp0_reg_6_ ( .D(n2604), .CK(clk), .Q(temp0[6]), .QN(n26587) );
  DFFXL temp0_reg_18_ ( .D(n2580), .CK(clk), .Q(temp0[18]), .QN(n26575) );
  DFFXL temp2_reg_4_ ( .D(n2609), .CK(clk), .Q(temp2[4]), .QN(n26540) );
  DFFXL temp0_reg_16_ ( .D(n2584), .CK(clk), .Q(temp0[16]), .QN(n26577) );
  DFFXL temp0_reg_5_ ( .D(n2606), .CK(clk), .Q(temp0[5]), .QN(n26588) );
  DFFXL temp2_reg_5_ ( .D(n2607), .CK(clk), .Q(temp2[5]), .QN(n26539) );
  DFFXL temp0_reg_17_ ( .D(n2582), .CK(clk), .Q(temp0[17]), .QN(n26576) );
  DFFXL temp0_reg_12_ ( .D(n2592), .CK(clk), .Q(temp0[12]), .QN(n26581) );
  DFFXL temp1_reg_16_ ( .D(n2538), .CK(clk), .Q(temp1[16]), .QN(n26554) );
  DFFXL temp1_reg_14_ ( .D(n2540), .CK(clk), .Q(temp1[14]), .QN(n26556) );
  DFFXL temp1_reg_13_ ( .D(n2541), .CK(clk), .Q(temp1[13]), .QN(n26557) );
  DFFXL temp1_reg_12_ ( .D(n2542), .CK(clk), .Q(temp1[12]), .QN(n26558) );
  DFFXL temp1_reg_9_ ( .D(n2545), .CK(clk), .Q(temp1[9]), .QN(n26561) );
  DFFXL temp1_reg_3_ ( .D(n2551), .CK(clk), .Q(temp1[3]), .QN(n26567) );
  DFFXL temp0_reg_15_ ( .D(n2586), .CK(clk), .Q(temp0[15]), .QN(n26578) );
  DFFXL temp0_reg_11_ ( .D(n2594), .CK(clk), .Q(temp0[11]), .QN(n26582) );
  DFFXL temp0_reg_14_ ( .D(n2588), .CK(clk), .Q(temp0[14]), .QN(n26579) );
  DFFXL temp0_reg_3_ ( .D(n2610), .CK(clk), .Q(temp0[3]), .QN(n26590) );
  DFFXL temp0_reg_8_ ( .D(n2600), .CK(clk), .Q(temp0[8]), .QN(n26585) );
  DFFXL temp2_reg_14_ ( .D(n2589), .CK(clk), .Q(temp2[14]), .QN(n26528) );
  DFFXL temp2_reg_18_ ( .D(n2581), .CK(clk), .Q(temp2[18]), .QN(n26524) );
  DFFXL temp2_reg_9_ ( .D(n2599), .CK(clk), .Q(temp2[9]), .QN(n26533) );
  DFFXL temp2_reg_7_ ( .D(n2603), .CK(clk), .Q(temp2[7]), .QN(n26537) );
  DFFXL temp0_reg_19_ ( .D(n2578), .CK(clk), .Q(temp0[19]), .QN(n26574) );
  DFFXL temp3_reg_13_ ( .D(mul5_out[13]), .CK(clk), .Q(temp3[13]) );
  DFFXL temp3_reg_12_ ( .D(mul5_out[12]), .CK(clk), .Q(temp3[12]) );
  DFFXL temp3_reg_10_ ( .D(mul5_out[10]), .CK(clk), .Q(temp3[10]) );
  DFFXL temp1_reg_21_ ( .D(n2533), .CK(clk), .Q(temp1[21]), .QN(n26549) );
  DFFXL temp0_reg_10_ ( .D(n2596), .CK(clk), .Q(temp0[10]), .QN(n26583) );
  DFFXL temp0_reg_9_ ( .D(n2598), .CK(clk), .Q(temp0[9]), .QN(n26584) );
  DFFXL temp0_reg_7_ ( .D(n2602), .CK(clk), .Q(temp0[7]), .QN(n26586) );
  DFFXL temp1_reg_10_ ( .D(n2544), .CK(clk), .Q(temp1[10]), .QN(n26560) );
  DFFXL temp2_reg_29_ ( .D(n2559), .CK(clk), .Q(temp2[29]), .QN(n26499) );
  DFFXL temp2_reg_26_ ( .D(n2565), .CK(clk), .Q(temp2[26]), .QN(n26503) );
  DFFXL temp2_reg_24_ ( .D(n2569), .CK(clk), .Q(temp2[24]), .QN(n26501) );
  DFFXL temp1_reg_5_ ( .D(n2549), .CK(clk), .Q(temp1[5]), .QN(n26565) );
  DFFXL temp2_reg_21_ ( .D(n2575), .CK(clk), .Q(temp2[21]), .QN(n26521) );
  DFFXL temp2_reg_28_ ( .D(n2561), .CK(clk), .Q(temp2[28]), .QN(n26498) );
  DFFXL temp2_reg_27_ ( .D(n2563), .CK(clk), .Q(temp2[27]), .QN(n26504) );
  DFFXL temp2_reg_25_ ( .D(n2567), .CK(clk), .Q(temp2[25]), .QN(n26502) );
  DFFXL temp2_reg_22_ ( .D(n2573), .CK(clk), .Q(temp2[22]), .QN(n26520) );
  DFFXL temp3_reg_11_ ( .D(mul5_out[11]), .CK(clk), .Q(temp3[11]) );
  DFFXL temp3_reg_20_ ( .D(mul5_out[20]), .CK(clk), .Q(temp3[20]) );
  DFFXL temp3_reg_19_ ( .D(mul5_out[19]), .CK(clk), .Q(temp3[19]) );
  DFFXL temp3_reg_21_ ( .D(mul5_out[21]), .CK(clk), .Q(temp3[21]) );
  DFFXL temp1_reg_18_ ( .D(n2536), .CK(clk), .Q(temp1[18]), .QN(n26552) );
  DFFSX4 sigma10_reg_2_ ( .D(n2266), .CK(clk), .SN(rst_n), .Q(n25900) );
  DFFHQXL temp3_reg_31_ ( .D(mul5_out[31]), .CK(clk), .Q(temp3[31]) );
  DFFHQXL learning_rate_reg_10_ ( .D(n2641), .CK(clk), .Q(learning_rate[10])
         );
  DFFSX2 cs_reg_2_ ( .D(n2489), .CK(clk), .SN(rst_n), .Q(n25886), .QN(cs[2])
         );
  AOI21XL M5_U3_U1_UEN0_0_3_1 ( .A0(M5_U3_U1_enc_tree_0__2__20_), .A1(
        M5_U3_U1_or2_inv_0__24_), .B0(M5_U3_U1_enc_tree_0__2__28_), .Y(
        M5_U3_U1_enc_tree_0__3__24_) );
  AOI21XL M1_U3_U1_UEN0_0_1_4 ( .A0(M1_a_14_), .A1(M1_U3_U1_or2_inv_0__18_), 
        .B0(M1_a_12_), .Y(M1_U3_U1_enc_tree_0__1__18_) );
  AOI21XL M1_U4_U1_UEN0_0_1_5 ( .A0(M1_b_10_), .A1(n6210), .B0(M1_b_8_), .Y(
        M1_U4_U1_enc_tree_0__1__22_) );
  AOI21XL M0_U3_U1_UEN0_2_3_1 ( .A0(M0_U3_U1_enc_tree_2__2__20_), .A1(
        M0_U3_U1_or2_inv_2__24_), .B0(M0_U3_U1_enc_tree_2__2__28_), .Y(
        M0_U3_U1_enc_tree_2__3__24_) );
  AOI21XL M4_U3_U1_UEN0_0_1_7 ( .A0(M4_a_2_), .A1(M4_U3_U1_or2_inv_0__30_), 
        .B0(M4_a_0_), .Y(M4_U3_U1_enc_tree_0__1__30_) );
  AOI21XL M1_U3_U1_UEN0_0_1_7 ( .A0(M1_a_2_), .A1(n13100), .B0(n13049), .Y(
        M1_U3_U1_enc_tree_0__1__30_) );
  AOI21XL M1_U3_U1_UEN0_0_1_6 ( .A0(M1_a_6_), .A1(M1_U3_U1_or2_inv_0__26_), 
        .B0(n25865), .Y(M1_U3_U1_enc_tree_0__1__26_) );
  AOI21XL M0_U4_U1_UEN0_0_1_7 ( .A0(M0_b_2_), .A1(n7056), .B0(M0_b_0_), .Y(
        M0_U4_U1_enc_tree_0__1__30_) );
  AOI21XL M1_U3_U1_UEN0_0_1_2 ( .A0(M1_a_22_), .A1(M1_U3_U1_or2_inv_0__10_), 
        .B0(M1_a_20_), .Y(M1_U3_U1_enc_tree_0__1__10_) );
  AOI21XL M3_U4_U1_UEN0_0_1_5 ( .A0(M4_mult_x_15_n1680), .A1(n6162), .B0(
        M3_mult_x_15_n1682), .Y(M3_U4_U1_enc_tree_0__1__22_) );
  DFFHQX2 valid_reg_0_ ( .D(N40), .CK(clk), .Q(valid[0]) );
  DFFSX1 y12_reg_17_ ( .D(n2427), .CK(clk), .SN(rst_n), .Q(n25963), .QN(
        y12[17]) );
  DFFHQXL learning_rate_reg_3_ ( .D(n2648), .CK(clk), .Q(learning_rate[3]) );
  DFFHQXL valid_reg_2_ ( .D(N42), .CK(clk), .Q(valid[2]) );
  DFFHQXL valid_reg_1_ ( .D(N41), .CK(clk), .Q(valid[1]) );
  DFFHQXL temp1_reg_31_ ( .D(n2619), .CK(clk), .Q(temp1[31]) );
  DFFHQXL temp0_reg_31_ ( .D(n2555), .CK(clk), .Q(temp0[31]) );
  DFFHQXL temp2_reg_31_ ( .D(n2618), .CK(clk), .Q(temp2[31]) );
  DFFHQXL learning_rate_reg_30_ ( .D(n2621), .CK(clk), .Q(learning_rate[30])
         );
  DFFHQXL learning_rate_reg_29_ ( .D(n2622), .CK(clk), .Q(learning_rate[29])
         );
  DFFHQXL learning_rate_reg_28_ ( .D(n2623), .CK(clk), .Q(learning_rate[28])
         );
  DFFHQXL learning_rate_reg_27_ ( .D(n2624), .CK(clk), .Q(learning_rate[27])
         );
  DFFHQXL learning_rate_reg_26_ ( .D(n2625), .CK(clk), .Q(learning_rate[26])
         );
  DFFHQXL learning_rate_reg_25_ ( .D(n2626), .CK(clk), .Q(learning_rate[25])
         );
  DFFHQXL learning_rate_reg_24_ ( .D(n2627), .CK(clk), .Q(learning_rate[24])
         );
  DFFHQXL learning_rate_reg_23_ ( .D(n2628), .CK(clk), .Q(learning_rate[23])
         );
  DFFHQXL learning_rate_reg_18_ ( .D(n2633), .CK(clk), .Q(learning_rate[18])
         );
  DFFHQXL learning_rate_reg_17_ ( .D(n2634), .CK(clk), .Q(learning_rate[17])
         );
  DFFHQXL learning_rate_reg_13_ ( .D(n2638), .CK(clk), .Q(learning_rate[13])
         );
  DFFHQXL learning_rate_reg_12_ ( .D(n2639), .CK(clk), .Q(learning_rate[12])
         );
  DFFHQXL learning_rate_reg_9_ ( .D(n2642), .CK(clk), .Q(learning_rate[9]) );
  DFFHQXL learning_rate_reg_8_ ( .D(n2643), .CK(clk), .Q(learning_rate[8]) );
  DFFHQXL learning_rate_reg_7_ ( .D(n2644), .CK(clk), .Q(learning_rate[7]) );
  DFFHQXL learning_rate_reg_5_ ( .D(n2646), .CK(clk), .Q(learning_rate[5]) );
  DFFHQXL learning_rate_reg_4_ ( .D(n2647), .CK(clk), .Q(learning_rate[4]) );
  DFFHQXL learning_rate_reg_2_ ( .D(n2649), .CK(clk), .Q(learning_rate[2]) );
  DFFHQXL learning_rate_reg_0_ ( .D(n2651), .CK(clk), .Q(learning_rate[0]) );
  DFFSX1 w1_reg_8__11_ ( .D(n2055), .CK(clk), .SN(rst_n), .QN(w1[267]) );
  AOI21XL M3_U4_U1_UEN0_0_3_1 ( .A0(M3_U4_U1_enc_tree_0__2__20_), .A1(
        M3_U4_U1_or2_inv_0__24_), .B0(M3_U4_U1_enc_tree_0__2__28_), .Y(
        M3_U4_U1_enc_tree_0__3__24_) );
  NOR2XL M4_U4_U1_UOR20_0_1_4 ( .A(M3_mult_x_15_b_15_), .B(M3_mult_x_15_b_13_), 
        .Y(M4_U4_U1_or2_tree_0__1__16_) );
  NAND2XL M2_U3_U1_UORT1_4_1 ( .A(M2_U3_U1_enc_tree_3__3__16_), .B(
        M2_U3_U1_enc_tree_3__3__24_), .Y(M2_U3_U1_enc_tree_4__4__16_) );
  NOR2XL M4_U4_U1_UORT0_3_3 ( .A(M4_U4_U1_enc_tree_2__2__24_), .B(
        M4_U4_U1_enc_tree_2__2__28_), .Y(M4_U4_U1_enc_tree_3__3__24_) );
  NOR2XL M4_U4_U1_UORT0_3_2 ( .A(M4_U4_U1_enc_tree_2__2__16_), .B(
        M4_U4_U1_enc_tree_2__2__20_), .Y(M4_U4_U1_enc_tree_3__3__16_) );
  NOR2XL M4_U3_U1_UORT0_3_2 ( .A(M4_U3_U1_enc_tree_2__2__16_), .B(
        M4_U3_U1_enc_tree_2__2__20_), .Y(M4_U3_U1_enc_tree_3__3__16_) );
  AOI21XL M1_U3_U1_UEN0_0_3_1 ( .A0(M1_U3_U1_enc_tree_0__2__20_), .A1(
        M1_U3_U1_or2_inv_0__24_), .B0(M1_U3_U1_enc_tree_0__2__28_), .Y(
        M1_U3_U1_enc_tree_0__3__24_) );
  AOI21XL M1_U4_U1_UEN0_0_3_1 ( .A0(M1_U4_U1_enc_tree_0__2__20_), .A1(
        M1_U4_U1_or2_inv_0__24_), .B0(M1_U4_U1_enc_tree_0__2__28_), .Y(
        M1_U4_U1_enc_tree_0__3__24_) );
  NOR2XL M1_U3_U1_UORT0_3_3 ( .A(M1_U3_U1_enc_tree_2__2__24_), .B(
        M1_U3_U1_enc_tree_2__2__28_), .Y(M1_U3_U1_enc_tree_3__3__24_) );
  NOR2XL M1_U3_U1_UORT0_3_2 ( .A(M1_U3_U1_enc_tree_2__2__16_), .B(
        M1_U3_U1_enc_tree_2__2__20_), .Y(M1_U3_U1_enc_tree_3__3__16_) );
  NOR2XL M1_U4_U1_UORT0_3_3 ( .A(M1_U4_U1_enc_tree_2__2__24_), .B(
        M1_U4_U1_enc_tree_2__2__28_), .Y(M1_U4_U1_enc_tree_3__3__24_) );
  NOR2XL M1_U4_U1_UORT0_3_2 ( .A(M1_U4_U1_enc_tree_2__2__16_), .B(
        M1_U4_U1_enc_tree_2__2__20_), .Y(M1_U4_U1_enc_tree_3__3__16_) );
  AOI21XL M2_U3_U1_UEN0_0_3_1 ( .A0(M2_U3_U1_enc_tree_0__2__20_), .A1(
        M2_U3_U1_or2_inv_0__24_), .B0(M2_U3_U1_enc_tree_0__2__28_), .Y(
        M2_U3_U1_enc_tree_0__3__24_) );
  AOI21XL M2_U3_U1_UEN0_1_3_1 ( .A0(M2_U3_U1_enc_tree_1__2__20_), .A1(
        M2_U3_U1_or2_inv_1__24_), .B0(M2_U3_U1_enc_tree_1__2__28_), .Y(
        M2_U3_U1_enc_tree_1__3__24_) );
  AOI21XL M2_U4_U1_UEN0_1_3_1 ( .A0(M2_U4_U1_enc_tree_1__2__20_), .A1(
        M2_U4_U1_or2_inv_1__24_), .B0(M2_U4_U1_enc_tree_1__2__28_), .Y(
        M2_U4_U1_enc_tree_1__3__24_) );
  NOR2XL M2_U4_U1_UORT0_3_3 ( .A(M2_U4_U1_enc_tree_2__2__24_), .B(
        M2_U4_U1_enc_tree_2__2__28_), .Y(M2_U4_U1_enc_tree_3__3__24_) );
  NOR2XL M2_U4_U1_UORT0_3_2 ( .A(M2_U4_U1_enc_tree_2__2__16_), .B(
        M2_U4_U1_enc_tree_2__2__20_), .Y(M2_U4_U1_enc_tree_3__3__16_) );
  NOR2XL M2_U3_U1_UORT0_3_3 ( .A(M2_U3_U1_enc_tree_2__2__24_), .B(
        M2_U3_U1_enc_tree_2__2__28_), .Y(M2_U3_U1_enc_tree_3__3__24_) );
  NOR2XL M2_U3_U1_UORT0_3_2 ( .A(M2_U3_U1_enc_tree_2__2__16_), .B(
        M2_U3_U1_enc_tree_2__2__20_), .Y(M2_U3_U1_enc_tree_3__3__16_) );
  AOI21XL M4_U3_U1_UEN0_1_3_1 ( .A0(M4_U3_U1_enc_tree_1__2__20_), .A1(
        M4_U3_U1_or2_inv_1__24_), .B0(M4_U3_U1_enc_tree_1__2__28_), .Y(
        M4_U3_U1_enc_tree_1__3__24_) );
  AOI21XL M3_U4_U1_UEN0_2_3_1 ( .A0(M4_U4_U1_enc_tree_2__2__20_), .A1(
        M3_U4_U1_or2_inv_2__24_), .B0(M4_U4_U1_enc_tree_2__2__28_), .Y(
        M3_U4_U1_enc_tree_2__3__24_) );
  AOI21XL M3_U4_U1_UEN0_1_3_1 ( .A0(M3_U4_U1_enc_tree_1__2__20_), .A1(
        M3_U4_U1_or2_inv_1__24_), .B0(M3_U4_U1_enc_tree_1__2__28_), .Y(
        M3_U4_U1_enc_tree_1__3__24_) );
  NAND2XL M4_U3_U1_UORT1_2_7 ( .A(M4_U3_U1_enc_tree_1__1__28_), .B(
        M4_U3_U1_enc_tree_1__1__30_), .Y(M4_U3_U1_enc_tree_2__2__28_) );
  NAND2XL M4_U3_U1_UORT1_2_6 ( .A(M4_U3_U1_enc_tree_1__1__24_), .B(
        M4_U3_U1_enc_tree_1__1__26_), .Y(M4_U3_U1_enc_tree_2__2__24_) );
  NAND2XL M4_U3_U1_UORT1_2_5 ( .A(M4_U3_U1_enc_tree_1__1__20_), .B(
        M4_U3_U1_enc_tree_1__1__22_), .Y(M4_U3_U1_enc_tree_2__2__20_) );
  NAND2XL M4_U3_U1_UORT1_2_4 ( .A(M4_U3_U1_enc_tree_1__1__16_), .B(
        M4_U3_U1_enc_tree_1__1__18_), .Y(M4_U3_U1_enc_tree_2__2__16_) );
  NOR2XL M5_U3_U1_UORT0_3_3 ( .A(M5_U3_U1_enc_tree_2__2__24_), .B(
        M5_U3_U1_enc_tree_2__2__28_), .Y(M5_U3_U1_enc_tree_3__3__24_) );
  NOR2XL M5_U3_U1_UORT0_3_2 ( .A(M5_U3_U1_enc_tree_2__2__16_), .B(
        M5_U3_U1_enc_tree_2__2__20_), .Y(M5_U3_U1_enc_tree_3__3__16_) );
  NOR2XL M3_U3_U1_UORT0_3_3 ( .A(M3_U3_U1_enc_tree_2__2__24_), .B(
        M3_U3_U1_enc_tree_2__2__28_), .Y(M3_U3_U1_enc_tree_3__3__24_) );
  NOR2XL M3_U3_U1_UORT0_3_2 ( .A(M3_U3_U1_enc_tree_2__2__16_), .B(
        M3_U3_U1_enc_tree_2__2__20_), .Y(M3_U3_U1_enc_tree_3__3__16_) );
  NOR2XL M0_U3_U1_UOR20_0_1_4 ( .A(n25869), .B(n23220), .Y(
        M0_U3_U1_or2_tree_0__1__16_) );
  NOR2XL M0_U4_U1_UOR20_0_1_4 ( .A(n25877), .B(n25878), .Y(
        M0_U4_U1_or2_tree_0__1__16_) );
  AOI21XL M0_U4_U1_UEN0_0_1_3 ( .A0(n25875), .A1(M0_U4_U1_or2_inv_0__14_), 
        .B0(n25876), .Y(M0_U4_U1_enc_tree_0__1__14_) );
  AOI21XL M0_U4_U1_UEN0_0_1_2 ( .A0(n25872), .A1(M0_U4_U1_or2_inv_0__10_), 
        .B0(n25873), .Y(M0_U4_U1_enc_tree_0__1__10_) );
  AOI21XL M0_U4_U1_UEN0_0_1_5 ( .A0(n25880), .A1(M0_U4_U1_or2_inv_0__22_), 
        .B0(n7475), .Y(M0_U4_U1_enc_tree_0__1__22_) );
  AOI21XL M0_U4_U1_UEN0_0_1_6 ( .A0(n25882), .A1(M0_U4_U1_or2_inv_0__26_), 
        .B0(M0_b_4_), .Y(M0_U4_U1_enc_tree_0__1__26_) );
  AOI21XL M0_U3_U1_UEN0_1_3_1 ( .A0(M0_U3_U1_enc_tree_1__2__20_), .A1(
        M0_U3_U1_or2_inv_1__24_), .B0(M0_U3_U1_enc_tree_1__2__28_), .Y(
        M0_U3_U1_enc_tree_1__3__24_) );
  AOI21XL M0_U4_U1_UEN0_1_3_1 ( .A0(M0_U4_U1_enc_tree_1__2__20_), .A1(
        M0_U4_U1_or2_inv_1__24_), .B0(M0_U4_U1_enc_tree_1__2__28_), .Y(
        M0_U4_U1_enc_tree_1__3__24_) );
  NOR2XL M0_U3_U1_UORT0_3_3 ( .A(M0_U3_U1_enc_tree_2__2__24_), .B(
        M0_U3_U1_enc_tree_2__2__28_), .Y(M0_U3_U1_enc_tree_3__3__24_) );
  NOR2XL M0_U3_U1_UORT0_3_2 ( .A(M0_U3_U1_enc_tree_2__2__16_), .B(
        M0_U3_U1_enc_tree_2__2__20_), .Y(M0_U3_U1_enc_tree_3__3__16_) );
  NOR2XL M0_U4_U1_UORT0_3_3 ( .A(M0_U4_U1_enc_tree_2__2__24_), .B(
        M0_U4_U1_enc_tree_2__2__28_), .Y(M0_U4_U1_enc_tree_3__3__24_) );
  NOR2XL M0_U4_U1_UORT0_3_2 ( .A(M0_U4_U1_enc_tree_2__2__16_), .B(
        M0_U4_U1_enc_tree_2__2__20_), .Y(M0_U4_U1_enc_tree_3__3__16_) );
  AOI21XL M0_U4_U1_UEN0_2_3_1 ( .A0(M0_U4_U1_enc_tree_2__2__20_), .A1(
        M0_U4_U1_or2_inv_2__24_), .B0(M0_U4_U1_enc_tree_2__2__28_), .Y(
        M0_U4_U1_enc_tree_2__3__24_) );
  AOI21XL M1_U3_U1_UEN0_2_3_1 ( .A0(M1_U3_U1_enc_tree_2__2__20_), .A1(
        M1_U3_U1_or2_inv_2__24_), .B0(M1_U3_U1_enc_tree_2__2__28_), .Y(
        M1_U3_U1_enc_tree_2__3__24_) );
  AOI21XL M1_U4_U1_UEN0_2_3_1 ( .A0(M1_U4_U1_enc_tree_2__2__20_), .A1(
        M1_U4_U1_or2_inv_2__24_), .B0(M1_U4_U1_enc_tree_2__2__28_), .Y(
        M1_U4_U1_enc_tree_2__3__24_) );
  AOI21XL M1_U4_U1_UEN0_1_3_1 ( .A0(M1_U4_U1_enc_tree_1__2__20_), .A1(
        M1_U4_U1_or2_inv_1__24_), .B0(M1_U4_U1_enc_tree_1__2__28_), .Y(
        M1_U4_U1_enc_tree_1__3__24_) );
  AOI21XL M1_U3_U1_UEN0_1_3_1 ( .A0(M1_U3_U1_enc_tree_1__2__20_), .A1(
        M1_U3_U1_or2_inv_1__24_), .B0(M1_U3_U1_enc_tree_1__2__28_), .Y(
        M1_U3_U1_enc_tree_1__3__24_) );
  AOI21XL M2_U3_U1_UEN0_2_3_1 ( .A0(M2_U3_U1_enc_tree_2__2__20_), .A1(
        M2_U3_U1_or2_inv_2__24_), .B0(M2_U3_U1_enc_tree_2__2__28_), .Y(
        M2_U3_U1_enc_tree_2__3__24_) );
  AOI21XL M2_U4_U1_UEN0_2_3_1 ( .A0(M2_U4_U1_enc_tree_2__2__20_), .A1(
        M2_U4_U1_or2_inv_2__24_), .B0(M2_U4_U1_enc_tree_2__2__28_), .Y(
        M2_U4_U1_enc_tree_2__3__24_) );
  AOI21XL M5_U3_U1_UEN0_2_3_1 ( .A0(M5_U3_U1_enc_tree_2__2__20_), .A1(
        M5_U3_U1_or2_inv_2__24_), .B0(M5_U3_U1_enc_tree_2__2__28_), .Y(
        M5_U3_U1_enc_tree_2__3__24_) );
  AOI21XL M5_U3_U1_UEN0_1_3_1 ( .A0(M5_U3_U1_enc_tree_1__2__20_), .A1(
        M5_U3_U1_or2_inv_1__24_), .B0(M5_U3_U1_enc_tree_1__2__28_), .Y(
        M5_U3_U1_enc_tree_1__3__24_) );
  AOI21XL M3_U3_U1_UEN0_2_3_1 ( .A0(M3_U3_U1_enc_tree_2__2__20_), .A1(
        M3_U3_U1_or2_inv_2__24_), .B0(M3_U3_U1_enc_tree_2__2__28_), .Y(
        M3_U3_U1_enc_tree_2__3__24_) );
  AOI21XL M3_U3_U1_UEN0_1_3_1 ( .A0(M3_U3_U1_enc_tree_1__2__20_), .A1(
        M3_U3_U1_or2_inv_1__24_), .B0(M3_U3_U1_enc_tree_1__2__28_), .Y(
        M3_U3_U1_enc_tree_1__3__24_) );
  AOI21XL M1_U3_U1_UEN0_0_1_3 ( .A0(n25864), .A1(M1_U3_U1_or2_inv_0__14_), 
        .B0(M1_a_16_), .Y(M1_U3_U1_enc_tree_0__1__14_) );
  NOR2XL M1_U4_U1_UOR20_0_1_5 ( .A(n25861), .B(n14030), .Y(
        M1_U4_U1_or2_tree_0__1__20_) );
  NOR2XL M1_U3_U1_UORT0_1_11 ( .A(n4567), .B(n4565), .Y(
        M1_U3_U1_enc_tree_1__1__22_) );
  AOI21XL M2_U4_U1_UEN0_0_1_7 ( .A0(M2_b_2_), .A1(n6076), .B0(M2_b_0_), .Y(
        M2_U4_U1_enc_tree_0__1__30_) );
  AOI21XL M4_U3_U1_UEN0_0_3_1 ( .A0(M4_U3_U1_enc_tree_0__2__20_), .A1(
        M4_U3_U1_or2_inv_0__24_), .B0(M4_U3_U1_enc_tree_0__2__28_), .Y(
        M4_U3_U1_enc_tree_0__3__24_) );
  NOR2XL M4_U3_U1_UORT0_3_3 ( .A(M4_U3_U1_enc_tree_2__2__24_), .B(
        M4_U3_U1_enc_tree_2__2__28_), .Y(M4_U3_U1_enc_tree_3__3__24_) );
  AOI21XL M3_U4_U1_UEN0_0_1_4 ( .A0(M3_mult_x_15_b_14_), .A1(
        M3_U4_U1_or2_inv_0__18_), .B0(n12561), .Y(M3_U4_U1_enc_tree_0__1__18_)
         );
  AOI21XL M3_U4_U1_UEN0_0_1_7 ( .A0(n12271), .A1(n5705), .B0(n2978), .Y(
        M3_U4_U1_enc_tree_0__1__30_) );
  AOI21XL M5_U3_U1_UEN0_0_1_5 ( .A0(M5_a_10_), .A1(n5729), .B0(M5_a_8_), .Y(
        M5_U3_U1_enc_tree_0__1__22_) );
  AOI21XL M5_U3_U1_UEN0_0_1_6 ( .A0(M5_a_6_), .A1(n16605), .B0(n4784), .Y(
        M5_U3_U1_enc_tree_0__1__26_) );
  AOI21XL M0_U3_U1_UEN0_0_3_1 ( .A0(M0_U3_U1_enc_tree_0__2__20_), .A1(
        M0_U3_U1_or2_inv_0__24_), .B0(M0_U3_U1_enc_tree_0__2__28_), .Y(
        M0_U3_U1_enc_tree_0__3__24_) );
  AOI21XL M0_U4_U1_UEN0_0_3_1 ( .A0(M0_U4_U1_enc_tree_0__2__20_), .A1(
        M0_U4_U1_or2_inv_0__24_), .B0(M0_U4_U1_enc_tree_0__2__28_), .Y(
        M0_U4_U1_enc_tree_0__3__24_) );
  AOI21XL M4_U3_U1_UEN0_2_3_1 ( .A0(M4_U3_U1_enc_tree_2__2__20_), .A1(
        M4_U3_U1_or2_inv_2__24_), .B0(M4_U3_U1_enc_tree_2__2__28_), .Y(
        M4_U3_U1_enc_tree_2__3__24_) );
  NAND2XL M4_U4_U1_UORT1_2_7 ( .A(M4_U4_U1_enc_tree_1__1__28_), .B(
        M4_U4_U1_enc_tree_1__1__30_), .Y(M4_U4_U1_enc_tree_2__2__28_) );
  NAND2XL M4_U4_U1_UORT1_2_6 ( .A(M4_U4_U1_enc_tree_1__1__24_), .B(
        M4_U4_U1_enc_tree_1__1__26_), .Y(M4_U4_U1_enc_tree_2__2__24_) );
  NAND2XL M4_U4_U1_UORT1_2_5 ( .A(M4_U4_U1_enc_tree_1__1__20_), .B(
        M4_U4_U1_enc_tree_1__1__22_), .Y(M4_U4_U1_enc_tree_2__2__20_) );
  NAND2XL M4_U4_U1_UORT1_2_4 ( .A(M4_U4_U1_enc_tree_1__1__16_), .B(
        M4_U4_U1_enc_tree_1__1__18_), .Y(M4_U4_U1_enc_tree_2__2__16_) );
  AOI21XL M3_U3_U1_UEN0_0_3_1 ( .A0(M3_U3_U1_enc_tree_0__2__20_), .A1(
        M3_U3_U1_or2_inv_0__24_), .B0(M3_U3_U1_enc_tree_0__2__28_), .Y(
        M3_U3_U1_enc_tree_0__3__24_) );
  AOI21XL M3_U3_U1_UEN0_0_1_2 ( .A0(M3_a_22_), .A1(n12751), .B0(M3_a_20_), .Y(
        M3_U3_U1_enc_tree_0__1__10_) );
  NAND2XL M1_U3_U1_UORT1_2_7 ( .A(M1_U3_U1_enc_tree_1__1__28_), .B(
        M1_U3_U1_enc_tree_1__1__30_), .Y(M1_U3_U1_enc_tree_2__2__28_) );
  NAND2XL M1_U3_U1_UORT1_2_6 ( .A(M1_U3_U1_enc_tree_1__1__24_), .B(
        M1_U3_U1_enc_tree_1__1__26_), .Y(M1_U3_U1_enc_tree_2__2__24_) );
  NAND2XL M1_U3_U1_UORT1_2_5 ( .A(M1_U3_U1_enc_tree_1__1__20_), .B(
        M1_U3_U1_enc_tree_1__1__22_), .Y(M1_U3_U1_enc_tree_2__2__20_) );
  NAND2XL M1_U3_U1_UORT1_2_4 ( .A(M1_U3_U1_enc_tree_1__1__16_), .B(
        M1_U3_U1_enc_tree_1__1__18_), .Y(M1_U3_U1_enc_tree_2__2__16_) );
  NAND2XL M1_U4_U1_UORT1_2_7 ( .A(M1_U4_U1_enc_tree_1__1__28_), .B(
        M1_U4_U1_enc_tree_1__1__30_), .Y(M1_U4_U1_enc_tree_2__2__28_) );
  NAND2XL M1_U4_U1_UORT1_2_6 ( .A(M1_U4_U1_enc_tree_1__1__24_), .B(
        M1_U4_U1_enc_tree_1__1__26_), .Y(M1_U4_U1_enc_tree_2__2__24_) );
  NAND2XL M1_U4_U1_UORT1_2_5 ( .A(M1_U4_U1_enc_tree_1__1__20_), .B(
        M1_U4_U1_enc_tree_1__1__22_), .Y(M1_U4_U1_enc_tree_2__2__20_) );
  NAND2XL M1_U4_U1_UORT1_2_4 ( .A(M1_U4_U1_enc_tree_1__1__16_), .B(
        M1_U4_U1_enc_tree_1__1__18_), .Y(M1_U4_U1_enc_tree_2__2__16_) );
  AOI21XL M2_U4_U1_UEN0_0_3_1 ( .A0(M2_U4_U1_enc_tree_0__2__20_), .A1(
        M2_U4_U1_or2_inv_0__24_), .B0(M2_U4_U1_enc_tree_0__2__28_), .Y(
        M2_U4_U1_enc_tree_0__3__24_) );
  NOR2XL M2_U4_U1_UOR20_0_1_4 ( .A(M2_b_15_), .B(M2_b_13_), .Y(
        M2_U4_U1_or2_tree_0__1__16_) );
  AOI21XL M2_U3_U1_UEN0_0_1_5 ( .A0(M2_a_10_), .A1(n9843), .B0(M2_a_8_), .Y(
        M2_U3_U1_enc_tree_0__1__22_) );
  NOR2XL M2_U3_U1_UOR20_0_1_6 ( .A(M2_a_7_), .B(M2_a_5_), .Y(
        M2_U3_U1_or2_tree_0__1__24_) );
  NAND2XL M2_U4_U1_UORT1_2_7 ( .A(M2_U4_U1_enc_tree_1__1__28_), .B(
        M2_U4_U1_enc_tree_1__1__30_), .Y(M2_U4_U1_enc_tree_2__2__28_) );
  NAND2XL M2_U4_U1_UORT1_2_6 ( .A(M2_U4_U1_enc_tree_1__1__24_), .B(
        M2_U4_U1_enc_tree_1__1__26_), .Y(M2_U4_U1_enc_tree_2__2__24_) );
  NAND2XL M2_U4_U1_UORT1_2_5 ( .A(M2_U4_U1_enc_tree_1__1__20_), .B(
        M2_U4_U1_enc_tree_1__1__22_), .Y(M2_U4_U1_enc_tree_2__2__20_) );
  NAND2XL M2_U4_U1_UORT1_2_4 ( .A(M2_U4_U1_enc_tree_1__1__16_), .B(
        M2_U4_U1_enc_tree_1__1__18_), .Y(M2_U4_U1_enc_tree_2__2__16_) );
  NAND2XL M2_U3_U1_UORT1_2_7 ( .A(M2_U3_U1_enc_tree_1__1__28_), .B(
        M2_U3_U1_enc_tree_1__1__30_), .Y(M2_U3_U1_enc_tree_2__2__28_) );
  NAND2XL M2_U3_U1_UORT1_2_6 ( .A(M2_U3_U1_enc_tree_1__1__24_), .B(
        M2_U3_U1_enc_tree_1__1__26_), .Y(M2_U3_U1_enc_tree_2__2__24_) );
  NAND2XL M2_U3_U1_UORT1_2_5 ( .A(M2_U3_U1_enc_tree_1__1__20_), .B(
        M2_U3_U1_enc_tree_1__1__22_), .Y(M2_U3_U1_enc_tree_2__2__20_) );
  NAND2XL M2_U3_U1_UORT1_2_4 ( .A(M2_U3_U1_enc_tree_1__1__16_), .B(
        M2_U3_U1_enc_tree_1__1__18_), .Y(M2_U3_U1_enc_tree_2__2__16_) );
  NOR2XL M4_U4_U1_UORT0_1_7 ( .A(n3201), .B(n11495), .Y(
        M4_U4_U1_enc_tree_1__1__14_) );
  NOR2XL M4_U4_U1_UORT0_1_6 ( .A(M3_mult_x_15_b_19_), .B(M5_b_18_), .Y(
        M4_U4_U1_enc_tree_1__1__12_) );
  NAND2XL M3_U4_U1_UOR21_1_2_3 ( .A(M4_U4_U1_enc_tree_1__1__24_), .B(
        M4_U4_U1_enc_tree_1__1__28_), .Y(M3_U4_U1_or2_tree_1__2__24_) );
  NAND2XL M3_U4_U1_UOR21_1_2_2 ( .A(M4_U4_U1_enc_tree_1__1__16_), .B(
        M4_U4_U1_enc_tree_1__1__20_), .Y(M3_U4_U1_or2_tree_1__2__16_) );
  NOR2XL M4_U4_U1_UORT0_1_5 ( .A(M3_mult_x_15_b_21_), .B(M3_mult_x_15_b_20_), 
        .Y(M4_U4_U1_enc_tree_1__1__10_) );
  NOR2XL M4_U4_U1_UORT0_1_12 ( .A(n3197), .B(M3_mult_x_15_b_6_), .Y(
        M4_U4_U1_enc_tree_1__1__24_) );
  NOR2XL M4_U4_U1_UORT0_1_8 ( .A(M3_mult_x_15_b_15_), .B(M3_mult_x_15_b_14_), 
        .Y(M4_U4_U1_enc_tree_1__1__16_) );
  NAND2XL M5_U3_U1_UORT1_2_7 ( .A(M5_U3_U1_enc_tree_1__1__28_), .B(
        M5_U3_U1_enc_tree_1__1__30_), .Y(M5_U3_U1_enc_tree_2__2__28_) );
  NAND2XL M5_U3_U1_UORT1_2_6 ( .A(M5_U3_U1_enc_tree_1__1__24_), .B(
        M5_U3_U1_enc_tree_1__1__26_), .Y(M5_U3_U1_enc_tree_2__2__24_) );
  NAND2XL M5_U3_U1_UORT1_2_5 ( .A(M5_U3_U1_enc_tree_1__1__20_), .B(
        M5_U3_U1_enc_tree_1__1__22_), .Y(M5_U3_U1_enc_tree_2__2__20_) );
  NAND2XL M5_U3_U1_UORT1_2_4 ( .A(M5_U3_U1_enc_tree_1__1__16_), .B(
        M5_U3_U1_enc_tree_1__1__18_), .Y(M5_U3_U1_enc_tree_2__2__16_) );
  NAND2XL M3_U3_U1_UORT1_2_7 ( .A(M3_U3_U1_enc_tree_1__1__28_), .B(
        M3_U3_U1_enc_tree_1__1__30_), .Y(M3_U3_U1_enc_tree_2__2__28_) );
  NAND2XL M3_U3_U1_UORT1_2_6 ( .A(M3_U3_U1_enc_tree_1__1__24_), .B(
        M3_U3_U1_enc_tree_1__1__26_), .Y(M3_U3_U1_enc_tree_2__2__24_) );
  NAND2XL M3_U3_U1_UORT1_2_5 ( .A(M3_U3_U1_enc_tree_1__1__20_), .B(
        M3_U3_U1_enc_tree_1__1__22_), .Y(M3_U3_U1_enc_tree_2__2__20_) );
  NAND2XL M3_U3_U1_UORT1_2_4 ( .A(M3_U3_U1_enc_tree_1__1__16_), .B(
        M3_U3_U1_enc_tree_1__1__18_), .Y(M3_U3_U1_enc_tree_2__2__16_) );
  NOR2XL M0_U3_U1_UOR20_0_1_5 ( .A(n25868), .B(n4789), .Y(
        M0_U3_U1_or2_tree_0__1__20_) );
  NOR2XL M0_U3_U1_UOR20_0_1_7 ( .A(n25866), .B(n21054), .Y(
        M0_U3_U1_or2_tree_0__1__28_) );
  NOR2XL M0_U4_U1_UOR20_0_1_5 ( .A(n25879), .B(M0_b_9_), .Y(
        M0_U4_U1_or2_tree_0__1__20_) );
  NAND2XL M0_U3_U1_UOR21_1_2_3 ( .A(M0_U3_U1_enc_tree_1__1__24_), .B(
        M0_U3_U1_enc_tree_1__1__28_), .Y(M0_U3_U1_or2_tree_1__2__24_) );
  NAND2XL M0_U4_U1_UOR21_1_2_3 ( .A(M0_U4_U1_enc_tree_1__1__24_), .B(
        M0_U4_U1_enc_tree_1__1__28_), .Y(M0_U4_U1_or2_tree_1__2__24_) );
  NAND2XL M0_U3_U1_UORT1_2_7 ( .A(M0_U3_U1_enc_tree_1__1__28_), .B(
        M0_U3_U1_enc_tree_1__1__30_), .Y(M0_U3_U1_enc_tree_2__2__28_) );
  NAND2XL M0_U3_U1_UORT1_2_6 ( .A(M0_U3_U1_enc_tree_1__1__24_), .B(
        M0_U3_U1_enc_tree_1__1__26_), .Y(M0_U3_U1_enc_tree_2__2__24_) );
  NAND2XL M0_U3_U1_UORT1_2_5 ( .A(M0_U3_U1_enc_tree_1__1__20_), .B(
        M0_U3_U1_enc_tree_1__1__22_), .Y(M0_U3_U1_enc_tree_2__2__20_) );
  NAND2XL M0_U3_U1_UORT1_2_4 ( .A(M0_U3_U1_enc_tree_1__1__16_), .B(
        M0_U3_U1_enc_tree_1__1__18_), .Y(M0_U3_U1_enc_tree_2__2__16_) );
  NAND2XL M0_U4_U1_UORT1_2_6 ( .A(M0_U4_U1_enc_tree_1__1__24_), .B(
        M0_U4_U1_enc_tree_1__1__26_), .Y(M0_U4_U1_enc_tree_2__2__24_) );
  NAND2XL M0_U4_U1_UORT1_2_7 ( .A(M0_U4_U1_enc_tree_1__1__28_), .B(
        M0_U4_U1_enc_tree_1__1__30_), .Y(M0_U4_U1_enc_tree_2__2__28_) );
  NAND2XL M0_U4_U1_UORT1_2_4 ( .A(M0_U4_U1_enc_tree_1__1__16_), .B(
        M0_U4_U1_enc_tree_1__1__18_), .Y(M0_U4_U1_enc_tree_2__2__16_) );
  NAND2XL M0_U4_U1_UORT1_2_5 ( .A(M0_U4_U1_enc_tree_1__1__20_), .B(
        M0_U4_U1_enc_tree_1__1__22_), .Y(M0_U4_U1_enc_tree_2__2__20_) );
  NOR2XL M0_U4_U1_UORT0_1_7 ( .A(M0_b_17_), .B(n25876), .Y(
        M0_U4_U1_enc_tree_1__1__14_) );
  NOR2XL M0_U4_U1_UORT0_1_6 ( .A(n25874), .B(n25875), .Y(
        M0_U4_U1_enc_tree_1__1__12_) );
  NOR2XL M1_U3_U1_UOR20_0_1_5 ( .A(M1_a_11_), .B(n4567), .Y(
        M1_U3_U1_or2_tree_0__1__20_) );
  NOR2XL M1_U3_U1_UORT0_1_7 ( .A(M1_a_17_), .B(M1_a_16_), .Y(
        M1_U3_U1_enc_tree_1__1__14_) );
  NOR2XL M1_U3_U1_UORT0_1_14 ( .A(M1_a_3_), .B(M1_a_2_), .Y(
        M1_U3_U1_enc_tree_1__1__28_) );
  NOR2XL M1_U3_U1_UORT0_1_13 ( .A(n13919), .B(M1_a_4_), .Y(
        M1_U3_U1_enc_tree_1__1__26_) );
  NOR2XL M1_U3_U1_UORT0_1_10 ( .A(M1_a_11_), .B(M1_a_10_), .Y(
        M1_U3_U1_enc_tree_1__1__20_) );
  NOR2XL M1_U3_U1_UORT0_1_9 ( .A(M1_a_13_), .B(M1_a_12_), .Y(
        M1_U3_U1_enc_tree_1__1__18_) );
  NOR2XL M1_U3_U1_UORT0_1_8 ( .A(M1_a_15_), .B(M1_a_14_), .Y(
        M1_U3_U1_enc_tree_1__1__16_) );
  NOR2XL M1_U4_U1_UORT0_1_13 ( .A(n4848), .B(M1_b_4_), .Y(
        M1_U4_U1_enc_tree_1__1__26_) );
  NOR2XL M1_U4_U1_UORT0_1_11 ( .A(n14030), .B(M1_b_8_), .Y(
        M1_U4_U1_enc_tree_1__1__22_) );
  NOR2XL M1_U4_U1_UORT0_1_10 ( .A(M1_b_11_), .B(M1_b_10_), .Y(
        M1_U4_U1_enc_tree_1__1__20_) );
  NOR2XL M1_U4_U1_UORT0_1_8 ( .A(M1_b_15_), .B(M1_b_14_), .Y(
        M1_U4_U1_enc_tree_1__1__16_) );
  NOR2XL M2_U4_U1_UORT0_1_7 ( .A(M2_b_17_), .B(n10335), .Y(
        M2_U4_U1_enc_tree_1__1__14_) );
  NOR2XL M2_U3_U1_UORT0_1_15 ( .A(M2_mult_x_15_a_1_), .B(M2_a_0_), .Y(
        M2_U3_U1_enc_tree_1__1__30_) );
  NOR2XL M2_U3_U1_UORT0_1_13 ( .A(M2_a_5_), .B(M2_a_4_), .Y(
        M2_U3_U1_enc_tree_1__1__26_) );
  NOR2XL M2_U3_U1_UORT0_1_14 ( .A(M2_a_3_), .B(M2_a_2_), .Y(
        M2_U3_U1_enc_tree_1__1__28_) );
  NOR2XL M2_U3_U1_UORT0_1_10 ( .A(n10324), .B(M2_a_10_), .Y(
        M2_U3_U1_enc_tree_1__1__20_) );
  NOR2XL M2_U3_U1_UORT0_1_12 ( .A(M2_a_7_), .B(M2_a_6_), .Y(
        M2_U3_U1_enc_tree_1__1__24_) );
  NOR2XL M2_U3_U1_UORT0_1_8 ( .A(M2_mult_x_15_n43), .B(M2_a_14_), .Y(
        M2_U3_U1_enc_tree_1__1__16_) );
  NOR2XL M2_U4_U1_UORT0_1_15 ( .A(n3182), .B(M2_b_0_), .Y(
        M2_U4_U1_enc_tree_1__1__30_) );
  NOR2XL M2_U4_U1_UORT0_1_9 ( .A(M2_b_13_), .B(M2_b_12_), .Y(
        M2_U4_U1_enc_tree_1__1__18_) );
  NOR2XL M2_U4_U1_UORT0_1_11 ( .A(n10311), .B(M2_b_8_), .Y(
        M2_U4_U1_enc_tree_1__1__22_) );
  NOR2XL M2_U4_U1_UORT0_1_12 ( .A(M2_b_7_), .B(M2_b_6_), .Y(
        M2_U4_U1_enc_tree_1__1__24_) );
  NAND2XL M5_U3_U1_UOR21_1_2_3 ( .A(M5_U3_U1_enc_tree_1__1__24_), .B(
        M5_U3_U1_enc_tree_1__1__28_), .Y(M5_U3_U1_or2_tree_1__2__24_) );
  NOR2XL M5_U3_U1_UORT0_1_12 ( .A(n4785), .B(M5_a_6_), .Y(
        M5_U3_U1_enc_tree_1__1__24_) );
  NOR2XL M5_U3_U1_UORT0_1_9 ( .A(n3199), .B(M5_a_12_), .Y(
        M5_U3_U1_enc_tree_1__1__18_) );
  NAND2XL M3_U3_U1_UOR21_1_2_3 ( .A(M3_U3_U1_enc_tree_1__1__24_), .B(
        M3_U3_U1_enc_tree_1__1__28_), .Y(M3_U3_U1_or2_tree_1__2__24_) );
  NOR2XL M3_U3_U1_UORT0_1_10 ( .A(M3_a_11_), .B(M3_a_10_), .Y(
        M3_U3_U1_enc_tree_1__1__20_) );
  NOR2XL M0_U3_U1_UORT0_1_14 ( .A(M0_a_3_), .B(M0_a_2_), .Y(
        M0_U3_U1_enc_tree_1__1__28_) );
  NOR2XL M0_U3_U1_UORT0_1_13 ( .A(n3209), .B(M0_a_4_), .Y(
        M0_U3_U1_enc_tree_1__1__26_) );
  NOR2XL M0_U3_U1_UORT0_1_11 ( .A(n4789), .B(M0_a_8_), .Y(
        M0_U3_U1_enc_tree_1__1__22_) );
  NOR2XL M0_U4_U1_UORT0_1_12 ( .A(M0_b_7_), .B(M0_b_6_), .Y(
        M0_U4_U1_enc_tree_1__1__24_) );
  NOR2XL M4_U4_U1_UOR20_0_1_6 ( .A(n3197), .B(n2974), .Y(
        M4_U4_U1_or2_tree_0__1__24_) );
  NAND2XL M3_U4_U1_UOR21_0_2_3 ( .A(M4_U4_U1_or2_tree_0__1__24_), .B(
        M4_U4_U1_or2_tree_0__1__28_), .Y(M3_U4_U1_or2_tree_0__2__24_) );
  NOR2XL M4_U4_U1_UOR20_0_1_5 ( .A(n3190), .B(M3_mult_x_15_b_9_), .Y(
        M4_U4_U1_or2_tree_0__1__20_) );
  NOR2XL M5_U3_U1_UOR20_0_1_6 ( .A(n4785), .B(n16614), .Y(
        M5_U3_U1_or2_tree_0__1__24_) );
  NAND2XL M5_U3_U1_UOR21_0_2_3 ( .A(M5_U3_U1_or2_tree_0__1__24_), .B(
        M5_U3_U1_or2_tree_0__1__28_), .Y(M5_U3_U1_or2_tree_0__2__24_) );
  NAND2XL M3_U3_U1_UOR21_0_2_3 ( .A(M3_U3_U1_or2_tree_0__1__24_), .B(
        M3_U3_U1_or2_tree_0__1__28_), .Y(M3_U3_U1_or2_tree_0__2__24_) );
  NAND2XL M2_U4_U1_UOR21_0_2_3 ( .A(M2_U4_U1_or2_tree_0__1__24_), .B(
        M2_U4_U1_or2_tree_0__1__28_), .Y(M2_U4_U1_or2_tree_0__2__24_) );
  NOR2XL M4_U4_U1_UORT0_1_15 ( .A(M3_mult_x_15_b_1_), .B(n3110), .Y(
        M4_U4_U1_enc_tree_1__1__30_) );
  NOR2XL M4_U4_U1_UORT0_1_14 ( .A(M3_mult_x_15_b_3_), .B(M3_mult_x_15_b_2_), 
        .Y(M4_U4_U1_enc_tree_1__1__28_) );
  NOR2XL M4_U4_U1_UORT0_1_13 ( .A(n2974), .B(n11499), .Y(
        M4_U4_U1_enc_tree_1__1__26_) );
  NOR2XL M4_U4_U1_UORT0_1_10 ( .A(M3_mult_x_15_b_11_), .B(n16884), .Y(
        M4_U4_U1_enc_tree_1__1__20_) );
  NOR2XL M4_U4_U1_UORT0_1_9 ( .A(M3_mult_x_15_b_13_), .B(n12561), .Y(
        M4_U4_U1_enc_tree_1__1__18_) );
  NOR2XL M4_U3_U1_UORT0_1_12 ( .A(n18118), .B(M4_a_6_), .Y(
        M4_U3_U1_enc_tree_1__1__24_) );
  NOR2XL M3_U3_U1_UOR20_0_1_7 ( .A(n11480), .B(n2980), .Y(
        M3_U3_U1_or2_tree_0__1__28_) );
  NAND2XL M0_U3_U1_UOR21_0_2_3 ( .A(M0_U3_U1_or2_tree_0__1__24_), .B(
        M0_U3_U1_or2_tree_0__1__28_), .Y(M0_U3_U1_or2_tree_0__2__24_) );
  NOR2XL M0_U4_U1_UOR20_0_1_6 ( .A(n25881), .B(M0_b_5_), .Y(
        M0_U4_U1_or2_tree_0__1__24_) );
  NAND2XL M0_U4_U1_UOR21_0_2_3 ( .A(M0_U4_U1_or2_tree_0__1__24_), .B(
        M0_U4_U1_or2_tree_0__1__28_), .Y(M0_U4_U1_or2_tree_0__2__24_) );
  NOR2XL M1_U4_U1_UORT0_1_6 ( .A(n25863), .B(M1_b_18_), .Y(
        M1_U4_U1_enc_tree_1__1__12_) );
  NOR2XL M1_U4_U1_UORT0_1_5 ( .A(n23173), .B(M1_b_20_), .Y(
        M1_U4_U1_enc_tree_1__1__10_) );
  NOR2XL M2_U3_U1_UORT0_1_6 ( .A(M2_a_19_), .B(M2_a_18_), .Y(
        M2_U3_U1_enc_tree_1__1__12_) );
  NOR2XL M2_U3_U1_UORT0_1_7 ( .A(n4808), .B(M2_a_16_), .Y(
        M2_U3_U1_enc_tree_1__1__14_) );
  NOR2XL M5_U3_U1_UORT0_1_15 ( .A(M5_mult_x_15_n1), .B(M5_a_0_), .Y(
        M5_U3_U1_enc_tree_1__1__30_) );
  NOR2XL M5_U3_U1_UORT0_1_14 ( .A(n3047), .B(M5_a_2_), .Y(
        M5_U3_U1_enc_tree_1__1__28_) );
  NOR2XL M5_U3_U1_UORT0_1_13 ( .A(n16614), .B(n4784), .Y(
        M5_U3_U1_enc_tree_1__1__26_) );
  NOR2XL M3_U3_U1_UORT0_1_15 ( .A(n2980), .B(n4776), .Y(
        M3_U3_U1_enc_tree_1__1__30_) );
  NOR2XL M0_U3_U1_UORT0_1_9 ( .A(n23220), .B(M0_a_12_), .Y(
        M0_U3_U1_enc_tree_1__1__18_) );
  NOR2XL M0_U4_U1_UORT0_1_10 ( .A(M0_b_11_), .B(M0_b_10_), .Y(
        M0_U4_U1_enc_tree_1__1__20_) );
  OR2XL M0_U4_U1_UOR20_0_1_3 ( .A(n25874), .B(M0_b_17_), .Y(
        M0_U4_U1_or2_tree_0__1__12_) );
  NOR2XL M4_U4_U1_UOR20_0_1_7 ( .A(n12279), .B(M3_mult_x_15_b_1_), .Y(
        M4_U4_U1_or2_tree_0__1__28_) );
  OR2XL M1_U3_U1_UOR20_0_1_3 ( .A(M1_a_19_), .B(M1_a_17_), .Y(
        M1_U3_U1_or2_tree_0__1__12_) );
  OR2XL M1_U4_U1_UOR20_0_1_3 ( .A(n25863), .B(n14228), .Y(
        M1_U4_U1_or2_tree_0__1__12_) );
  OR2XL M2_U3_U1_UOR20_0_1_3 ( .A(M2_a_19_), .B(n4808), .Y(
        M2_U3_U1_or2_tree_0__1__12_) );
  NOR2XL M2_U3_U1_UOR20_0_1_7 ( .A(n9904), .B(M2_mult_x_15_a_1_), .Y(
        M2_U3_U1_or2_tree_0__1__28_) );
  OR2XL M4_U4_U1_UOR20_0_1_3 ( .A(M3_mult_x_15_b_19_), .B(n3201), .Y(
        M4_U4_U1_or2_tree_0__1__12_) );
  DFFSX1 sigma10_reg_11_ ( .D(n2275), .CK(clk), .SN(rst_n), .Q(n26234), .QN(
        sigma10[11]) );
  DFFSX1 y10_reg_15_ ( .D(n2422), .CK(clk), .SN(rst_n), .Q(n26224), .QN(
        y10[15]) );
  DFFSX1 y10_reg_19_ ( .D(n2430), .CK(clk), .SN(rst_n), .Q(n26229), .QN(
        y10[19]) );
  DFFSX1 y10_reg_24_ ( .D(n2440), .CK(clk), .SN(rst_n), .Q(n26291), .QN(
        y10[24]) );
  DFFSX1 y12_reg_5_ ( .D(n2403), .CK(clk), .SN(rst_n), .Q(n25975), .QN(y12[5])
         );
  DFFSX1 y12_reg_15_ ( .D(n2423), .CK(clk), .SN(rst_n), .Q(n25965), .QN(
        y12[15]) );
  DFFRX1 y10_reg_28_ ( .D(n25859), .CK(clk), .RN(rst_n), .Q(y10[28]) );
  DFFXL temp2_reg_12_ ( .D(n2593), .CK(clk), .Q(temp2[12]), .QN(n26530) );
  DFFSX1 y11_reg_2_ ( .D(n2458), .CK(clk), .SN(rst_n), .Q(n25954), .QN(y11[2])
         );
  DFFSX1 y11_reg_26_ ( .D(n2482), .CK(clk), .SN(rst_n), .Q(n26185), .QN(
        y11[26]) );
  DFFSX1 w2_reg_1__14_ ( .D(n2182), .CK(clk), .SN(rst_n), .Q(n26436), .QN(
        w2[46]) );
  DFFSX1 y12_reg_29_ ( .D(n2451), .CK(clk), .SN(rst_n), .Q(n26188), .QN(
        y12[29]) );
  DFFSX1 y11_reg_28_ ( .D(n2484), .CK(clk), .SN(rst_n), .Q(n26186), .QN(
        y11[28]) );
  DFFSX1 y11_reg_24_ ( .D(n2480), .CK(clk), .SN(rst_n), .Q(n26187), .QN(
        y11[24]) );
  DFFSX1 y11_reg_25_ ( .D(n2481), .CK(clk), .SN(rst_n), .Q(n25936), .QN(
        y11[25]) );
  DFFSX1 y11_reg_27_ ( .D(n2483), .CK(clk), .SN(rst_n), .Q(n25937), .QN(
        y11[27]) );
  DFFSX1 y11_reg_29_ ( .D(n2485), .CK(clk), .SN(rst_n), .Q(n25935), .QN(
        y11[29]) );
  DFFSX1 y11_reg_9_ ( .D(n2465), .CK(clk), .SN(rst_n), .Q(n25891), .QN(y11[9])
         );
  DFFSX1 y11_reg_23_ ( .D(n2479), .CK(clk), .SN(rst_n), .Q(n26142), .QN(
        y11[23]) );
  DFFSX1 y11_reg_6_ ( .D(n2462), .CK(clk), .SN(rst_n), .Q(n25950), .QN(y11[6])
         );
  DFFSX1 w2_reg_2__22_ ( .D(n2222), .CK(clk), .SN(rst_n), .QN(w2[86]) );
  DFFSX1 y11_reg_30_ ( .D(n2486), .CK(clk), .SN(rst_n), .Q(n25957), .QN(
        y11[30]) );
  DFFSX1 y12_reg_28_ ( .D(n2449), .CK(clk), .SN(rst_n), .Q(n26191), .QN(
        y12[28]) );
  DFFSX1 y12_reg_24_ ( .D(n2441), .CK(clk), .SN(rst_n), .Q(n26193), .QN(
        y12[24]) );
  DFFSX1 y12_reg_26_ ( .D(n2445), .CK(clk), .SN(rst_n), .Q(n26194), .QN(
        y12[26]) );
  DFFSX1 y12_reg_27_ ( .D(n2447), .CK(clk), .SN(rst_n), .Q(n26190), .QN(
        y12[27]) );
  DFFSX1 y12_reg_16_ ( .D(n2425), .CK(clk), .SN(rst_n), .Q(n25964), .QN(
        y12[16]) );
  DFFSX1 y12_reg_12_ ( .D(n2417), .CK(clk), .SN(rst_n), .Q(n25968), .QN(
        y12[12]) );
  DFFSX1 y12_reg_2_ ( .D(n2397), .CK(clk), .SN(rst_n), .Q(n25978), .QN(y12[2])
         );
  DFFSX1 y12_reg_4_ ( .D(n2401), .CK(clk), .SN(rst_n), .Q(n25976), .QN(y12[4])
         );
  DFFSX1 y12_reg_6_ ( .D(n2405), .CK(clk), .SN(rst_n), .Q(n25974), .QN(y12[6])
         );
  DFFSX1 y12_reg_19_ ( .D(n2431), .CK(clk), .SN(rst_n), .Q(n25961), .QN(
        y12[19]) );
  DFFSX1 y12_reg_13_ ( .D(n2419), .CK(clk), .SN(rst_n), .Q(n25967), .QN(
        y12[13]) );
  DFFSX1 y12_reg_11_ ( .D(n2415), .CK(clk), .SN(rst_n), .Q(n25969), .QN(
        y12[11]) );
  DFFSX1 y12_reg_10_ ( .D(n2413), .CK(clk), .SN(rst_n), .Q(n25970), .QN(
        y12[10]) );
  DFFSX1 y12_reg_1_ ( .D(n2395), .CK(clk), .SN(rst_n), .Q(n25979), .QN(y12[1])
         );
  DFFSX1 y12_reg_9_ ( .D(n2411), .CK(clk), .SN(rst_n), .Q(n25971), .QN(y12[9])
         );
  DFFSX1 y12_reg_25_ ( .D(n2443), .CK(clk), .SN(rst_n), .Q(n26189), .QN(
        y12[25]) );
  DFFSX1 w2_reg_0__8_ ( .D(n2144), .CK(clk), .SN(rst_n), .Q(n26003), .QN(w2[8]) );
  DFFSX1 y10_reg_27_ ( .D(n2446), .CK(clk), .SN(rst_n), .Q(n26299), .QN(
        y10[27]) );
  DFFSX1 y10_reg_2_ ( .D(n2396), .CK(clk), .SN(rst_n), .Q(n25896), .QN(y10[2])
         );
  DFFSX1 y10_reg_0_ ( .D(n2392), .CK(clk), .SN(rst_n), .Q(n26226), .QN(y10[0])
         );
  DFFSX1 y10_reg_1_ ( .D(n2394), .CK(clk), .SN(rst_n), .Q(n25895), .QN(y10[1])
         );
  DFFSX1 y10_reg_8_ ( .D(n2408), .CK(clk), .SN(rst_n), .Q(n26220), .QN(y10[8])
         );
  DFFSX1 y20_reg_21_ ( .D(n2381), .CK(clk), .SN(rst_n), .Q(n26167), .QN(
        y20[21]) );
  DFFSX1 y10_reg_25_ ( .D(n2442), .CK(clk), .SN(rst_n), .Q(n26289), .QN(
        y10[25]) );
  DFFSX1 y10_reg_17_ ( .D(n2426), .CK(clk), .SN(rst_n), .Q(n26228), .QN(
        y10[17]) );
  DFFSX1 y10_reg_18_ ( .D(n2428), .CK(clk), .SN(rst_n), .Q(n25993), .QN(
        y10[18]) );
  DFFSX1 y10_reg_5_ ( .D(n2402), .CK(clk), .SN(rst_n), .Q(n26217), .QN(y10[5])
         );
  DFFSX1 y10_reg_22_ ( .D(n2436), .CK(clk), .SN(rst_n), .Q(n26231), .QN(
        y10[22]) );
  DFFSX1 y10_reg_6_ ( .D(n2404), .CK(clk), .SN(rst_n), .Q(n26218), .QN(y10[6])
         );
  DFFSX1 y10_reg_20_ ( .D(n2432), .CK(clk), .SN(rst_n), .Q(n26230), .QN(
        y10[20]) );
  DFFSX1 y10_reg_14_ ( .D(n2420), .CK(clk), .SN(rst_n), .Q(n26223), .QN(
        y10[14]) );
  DFFSX1 y10_reg_12_ ( .D(n2416), .CK(clk), .SN(rst_n), .Q(n26221), .QN(
        y10[12]) );
  DFFSX1 y20_reg_5_ ( .D(n2365), .CK(clk), .SN(rst_n), .Q(n26183), .QN(y20[5])
         );
  DFFSX1 y20_reg_12_ ( .D(n2372), .CK(clk), .SN(rst_n), .Q(n26177), .QN(
        y20[12]) );
  DFFSX1 y20_reg_14_ ( .D(n2374), .CK(clk), .SN(rst_n), .Q(n26175), .QN(
        y20[14]) );
  DFFSX1 y20_reg_4_ ( .D(n2364), .CK(clk), .SN(rst_n), .Q(n26184), .QN(y20[4])
         );
  DFFSX1 sigma10_reg_23_ ( .D(n2287), .CK(clk), .SN(rst_n), .Q(n26286), .QN(
        sigma10[23]) );
  DFFSX1 sigma10_reg_24_ ( .D(n2288), .CK(clk), .SN(rst_n), .Q(n26282), .QN(
        sigma10[24]) );
  DFFSX1 sigma10_reg_26_ ( .D(n2290), .CK(clk), .SN(rst_n), .Q(n26297), .QN(
        sigma10[26]) );
  DFFSX1 sigma10_reg_25_ ( .D(n2289), .CK(clk), .SN(rst_n), .Q(n26411), .QN(
        sigma10[25]) );
  DFFSX1 sigma12_reg_23_ ( .D(n2342), .CK(clk), .SN(rst_n), .Q(n26453), .QN(
        sigma12[23]) );
  DFFSX1 sigma12_reg_24_ ( .D(n2344), .CK(clk), .SN(rst_n), .Q(n26137), .QN(
        sigma12[24]) );
  DFFSX1 sigma10_reg_27_ ( .D(n2291), .CK(clk), .SN(rst_n), .Q(n26410), .QN(
        sigma10[27]) );
  DFFSX1 sigma10_reg_28_ ( .D(n2292), .CK(clk), .SN(rst_n), .Q(n26302), .QN(
        sigma10[28]) );
  DFFSX1 sigma12_reg_25_ ( .D(n2346), .CK(clk), .SN(rst_n), .Q(n26414), .QN(
        sigma12[25]) );
  DFFSX1 sigma10_reg_30_ ( .D(n2294), .CK(clk), .SN(rst_n), .Q(n26303), .QN(
        sigma10[30]) );
  DFFSX1 sigma10_reg_29_ ( .D(n2293), .CK(clk), .SN(rst_n), .Q(n26412), .QN(
        sigma10[29]) );
  DFFSX1 sigma12_reg_29_ ( .D(n2354), .CK(clk), .SN(rst_n), .Q(n26415), .QN(
        sigma12[29]) );
  DFFSX2 o_valid_reg ( .D(n26595), .CK(clk), .SN(rst_n), .Q(n26487), .QN(n2972) );
  OAI2BB1XL U3297 ( .A0N(n21167), .A1N(n24248), .B0(n4837), .Y(n2336) );
  OAI2BB1X1 U3298 ( .A0N(n25767), .A1N(n25293), .B0(n4839), .Y(n2298) );
  OAI2BB1X1 U3299 ( .A0N(n25767), .A1N(n24116), .B0(n4838), .Y(n2300) );
  OAI21XL U3300 ( .A0(n24656), .A1(n3059), .B0(n24653), .Y(n24654) );
  INVX1 U3301 ( .A(n24264), .Y(mul5_out[0]) );
  OAI21XL U3302 ( .A0(n25506), .A1(n3059), .B0(n3818), .Y(n3819) );
  OAI21XL U3303 ( .A0(n24616), .A1(n3059), .B0(n24613), .Y(n24614) );
  INVXL U3304 ( .A(n23604), .Y(n23721) );
  OAI21XL U3305 ( .A0(n24843), .A1(n24632), .B0(n24840), .Y(n24841) );
  OAI21XL U3306 ( .A0(n24868), .A1(n3024), .B0(n24865), .Y(n24866) );
  OAI21XL U3307 ( .A0(n25594), .A1(n3024), .B0(n24499), .Y(n24500) );
  OAI21XL U3308 ( .A0(n24697), .A1(n3024), .B0(n24694), .Y(n24695) );
  OAI21XL U3309 ( .A0(n24515), .A1(n3024), .B0(n20998), .Y(n20999) );
  OAI21XL U3310 ( .A0(n4081), .A1(n4875), .B0(n24175), .Y(n5043) );
  OAI21XL U3311 ( .A0(n25176), .A1(n3111), .B0(n25175), .Y(n25177) );
  OAI2BB1X1 U3312 ( .A0N(n3136), .A1N(n20943), .B0(n5850), .Y(mul5_out[17]) );
  OAI21XL U3313 ( .A0(n25758), .A1(n25757), .B0(n25756), .Y(n25759) );
  OAI21XL U3314 ( .A0(n25093), .A1(n3024), .B0(n25091), .Y(n25092) );
  OAI21XL U3315 ( .A0(n25842), .A1(n3024), .B0(n25672), .Y(n25673) );
  OAI21XL U3316 ( .A0(n25722), .A1(n3024), .B0(n24415), .Y(n24416) );
  OAI2BB1X1 U3317 ( .A0N(n3136), .A1N(n21049), .B0(n3630), .Y(mul5_out[19]) );
  OAI2BB1X1 U3318 ( .A0N(n5336), .A1N(n21049), .B0(n4167), .Y(mul5_out[18]) );
  OAI2BB1X1 U3319 ( .A0N(n3136), .A1N(n20343), .B0(n6044), .Y(mul5_out[5]) );
  OAI2BB1X1 U3320 ( .A0N(n20747), .A1N(n3136), .B0(n20344), .Y(mul5_out[4]) );
  OAI2BB1X1 U3321 ( .A0N(n20337), .A1N(n3136), .B0(n17449), .Y(mul5_out[9]) );
  OAI2BB1X1 U3322 ( .A0N(n20742), .A1N(n3136), .B0(n20338), .Y(mul5_out[8]) );
  OAI21XL U3323 ( .A0(n25197), .A1(n3111), .B0(n25196), .Y(n25198) );
  OAI21XL U3324 ( .A0(n24256), .A1(n24119), .B0(n24118), .Y(n24120) );
  OAI21XL U3325 ( .A0(n24256), .A1(n24142), .B0(n24141), .Y(n24143) );
  OAI21XL U3326 ( .A0(n24256), .A1(n24165), .B0(n24164), .Y(n24166) );
  OAI21XL U3327 ( .A0(n24256), .A1(n24255), .B0(n24254), .Y(n24258) );
  OAI21XL U3328 ( .A0(n24132), .A1(n3111), .B0(n24131), .Y(n24133) );
  AOI2BB1X1 U3329 ( .A0N(n24656), .A1N(n4582), .B0(n5916), .Y(n5915) );
  AOI2BB1X1 U3330 ( .A0N(n24984), .A1N(n4586), .B0(n6006), .Y(n6005) );
  AOI2BB1X1 U3331 ( .A0N(n24936), .A1N(n4584), .B0(n5965), .Y(n5341) );
  AOI22X1 U3332 ( .A0(n3131), .A1(n5366), .B0(n3467), .B1(n24140), .Y(n21029)
         );
  AOI2BB1X1 U3333 ( .A0N(n24888), .A1N(n4581), .B0(n4810), .Y(n4857) );
  AOI2BB1X1 U3334 ( .A0N(n23593), .A1N(n4583), .B0(n3531), .Y(n3530) );
  AOI2BB1X1 U3335 ( .A0N(n23912), .A1N(n4583), .B0(n23911), .Y(n23913) );
  AOI2BB1X1 U3336 ( .A0N(n23825), .A1N(n4583), .B0(n5597), .Y(n3515) );
  OAI21X1 U3337 ( .A0(n5710), .A1(n5695), .B0(n5694), .Y(mul5_out[22]) );
  NOR2X2 U3338 ( .A(n4342), .B(n3121), .Y(n25636) );
  OAI2BB1X1 U3339 ( .A0N(n23620), .A1N(n3455), .B0(n4546), .Y(n25740) );
  OAI2BB1X1 U3340 ( .A0N(n20882), .A1N(n3455), .B0(n4555), .Y(n23701) );
  INVXL U3341 ( .A(n24319), .Y(n24315) );
  OAI2BB1X1 U3342 ( .A0N(n3081), .A1N(n23435), .B0(n4264), .Y(n24655) );
  AOI22X1 U3343 ( .A0(n3128), .A1(n20754), .B0(n23522), .B1(n23534), .Y(n24735) );
  AOI22X1 U3344 ( .A0(n23724), .A1(n19104), .B0(n3128), .B1(n23462), .Y(n24515) );
  NAND2X1 U3345 ( .A(n20939), .B(n3136), .Y(n5694) );
  AOI22X1 U3346 ( .A0(n3128), .A1(n23944), .B0(n23926), .B1(n19104), .Y(n24616) );
  NAND2X1 U3347 ( .A(n20933), .B(n5336), .Y(n3630) );
  AOI22X1 U3348 ( .A0(n3128), .A1(n23536), .B0(n23535), .B1(n23534), .Y(n24843) );
  OAI2BB1X2 U3349 ( .A0N(n3455), .A1N(n23894), .B0(n3580), .Y(n24743) );
  AOI22X1 U3350 ( .A0(n20814), .A1(n19104), .B0(n23535), .B1(n3128), .Y(n24821) );
  AOI22X1 U3351 ( .A0(n23522), .A1(n3128), .B0(n19104), .B1(n23521), .Y(n24697) );
  NAND2X1 U3352 ( .A(n3136), .B(n20936), .Y(n3950) );
  AOI22X1 U3353 ( .A0(n23724), .A1(n3128), .B0(n23723), .B1(n23722), .Y(n25594) );
  AOI22X1 U3354 ( .A0(n23944), .A1(n19104), .B0(n3128), .B1(n23945), .Y(n25506) );
  OAI2BB1X2 U3355 ( .A0N(n3139), .A1N(n23806), .B0(n20621), .Y(n3602) );
  AOI22X1 U3356 ( .A0(n23626), .A1(n4267), .B0(n23627), .B1(n3081), .Y(n24491)
         );
  NAND2XL U3357 ( .A(n20733), .B(n5336), .Y(n5721) );
  AOI22X1 U3358 ( .A0(n23925), .A1(n3128), .B0(n3325), .B1(n19104), .Y(n24582)
         );
  XNOR2XL U3359 ( .A(n3357), .B(n20692), .Y(n21051) );
  NAND2X1 U3360 ( .A(n3548), .B(n3547), .Y(n25733) );
  NAND2X1 U3361 ( .A(n3576), .B(n3575), .Y(n23758) );
  NAND2XL U3362 ( .A(n3491), .B(n3490), .Y(n24526) );
  NAND2XL U3363 ( .A(n3493), .B(n3492), .Y(n25738) );
  AOI22X1 U3364 ( .A0(n20620), .A1(n3139), .B0(n3455), .B1(n23612), .Y(n23825)
         );
  AOI22X2 U3365 ( .A0(n20716), .A1(n3128), .B0(n20712), .B1(n23722), .Y(n25731) );
  AOI22X1 U3366 ( .A0(n3001), .A1(n5336), .B0(n20733), .B1(n3136), .Y(n24200)
         );
  AOI22X1 U3367 ( .A0(n25553), .A1(n4215), .B0(n4220), .B1(n23479), .Y(n24132)
         );
  AOI21XL U3368 ( .A0(n4215), .A1(n25591), .B0(n4256), .Y(n24115) );
  AOI22X1 U3369 ( .A0(n3353), .A1(n4382), .B0(n17458), .B1(n3131), .Y(n20691)
         );
  NAND2XL U3370 ( .A(n4295), .B(n4291), .Y(n24535) );
  OAI2BB1X1 U3371 ( .A0N(n3455), .A1N(n23619), .B0(n3502), .Y(n24548) );
  NAND3BXL U3372 ( .AN(n3004), .B(n4498), .C(n4497), .Y(n25679) );
  NOR2X1 U3373 ( .A(n3772), .B(n3770), .Y(n25197) );
  AOI21X1 U3374 ( .A0(n20792), .A1(n5229), .B0(n5230), .Y(n25709) );
  AOI2BB1X1 U3375 ( .A0N(n24631), .A1N(n3227), .B0(n3820), .Y(n3818) );
  AOI211X1 U3376 ( .A0(n20778), .A1(n5911), .B0(n20777), .C0(n25127), .Y(
        n25176) );
  CLKINVX3 U3377 ( .A(n23235), .Y(n23257) );
  BUFX4 U3378 ( .A(n24617), .Y(n3029) );
  INVX1 U3379 ( .A(n3139), .Y(n5589) );
  OAI21XL U3380 ( .A0(n20789), .A1(n4369), .B0(n24380), .Y(n5230) );
  XOR2X1 U3381 ( .A(n5515), .B(n23548), .Y(n24206) );
  XOR2X1 U3382 ( .A(n5880), .B(n19021), .Y(n24210) );
  XOR2X1 U3383 ( .A(n5025), .B(n14689), .Y(n23703) );
  OAI21XL U3384 ( .A0(n24439), .A1(n24095), .B0(n24094), .Y(n25227) );
  OAI21XL U3385 ( .A0(n24439), .A1(n24344), .B0(n24343), .Y(n24373) );
  OAI21XL U3386 ( .A0(n24439), .A1(n24303), .B0(n24302), .Y(n25816) );
  OAI21XL U3387 ( .A0(n24439), .A1(n24438), .B0(n24437), .Y(n25671) );
  OAI21XL U3388 ( .A0(n24439), .A1(n24312), .B0(n24311), .Y(n25810) );
  OAI21XL U3389 ( .A0(n24439), .A1(n24298), .B0(n24297), .Y(n25090) );
  XOR2X1 U3390 ( .A(n20992), .B(n4442), .Y(n23724) );
  NAND2X1 U3391 ( .A(n20847), .B(n3139), .Y(n3580) );
  NAND2X1 U3392 ( .A(n3139), .B(n23620), .Y(n3502) );
  XOR2X1 U3393 ( .A(n4010), .B(n20669), .Y(n24237) );
  XOR2X1 U3394 ( .A(n17490), .B(n20270), .Y(n23536) );
  NAND2XL U3395 ( .A(n20900), .B(n3139), .Y(n6025) );
  XNOR2X1 U3396 ( .A(n20325), .B(n20324), .Y(n5366) );
  NAND2XL U3397 ( .A(n23612), .B(n3139), .Y(n3548) );
  NAND2X1 U3398 ( .A(n4267), .B(n23627), .Y(n5153) );
  NAND2XL U3399 ( .A(n3455), .B(n23611), .Y(n3547) );
  NAND2XL U3400 ( .A(n3455), .B(n20819), .Y(n3576) );
  NAND2XL U3401 ( .A(n3139), .B(n23619), .Y(n3491) );
  XOR2X1 U3402 ( .A(n5665), .B(n20355), .Y(n20733) );
  XOR2X1 U3403 ( .A(n5799), .B(n19050), .Y(n24199) );
  NAND2XL U3404 ( .A(n3483), .B(n3139), .Y(n3489) );
  NAND2XL U3405 ( .A(n24135), .B(n3131), .Y(n3468) );
  XOR2X1 U3406 ( .A(n23735), .B(n3147), .Y(n25502) );
  XOR2XL U3407 ( .A(n20664), .B(n20663), .Y(n5340) );
  XOR2X1 U3408 ( .A(n4214), .B(n23530), .Y(n25552) );
  NAND2X1 U3409 ( .A(n4000), .B(n3131), .Y(n3999) );
  NAND2X1 U3410 ( .A(n3976), .B(n3353), .Y(n5953) );
  XOR2XL U3411 ( .A(n20976), .B(n23444), .Y(n23879) );
  XNOR2X1 U3412 ( .A(n19102), .B(n5191), .Y(n23741) );
  XOR2X1 U3413 ( .A(n5386), .B(n5385), .Y(n4283) );
  NAND3BX1 U3414 ( .AN(n5426), .B(n5425), .C(n3409), .Y(n25378) );
  NAND3X1 U3415 ( .A(n5383), .B(n5382), .C(n5381), .Y(n23747) );
  XNOR2X1 U3416 ( .A(n23740), .B(n5749), .Y(n23945) );
  NAND2X1 U3417 ( .A(n5271), .B(n5266), .Y(n24696) );
  XOR2X1 U3418 ( .A(n5822), .B(n23455), .Y(n25591) );
  XOR2X1 U3419 ( .A(n4887), .B(n4886), .Y(n24236) );
  NAND3X1 U3420 ( .A(n6022), .B(n6132), .C(n6031), .Y(n24397) );
  OAI21X1 U3421 ( .A0(n4190), .A1(n5914), .B0(n5913), .Y(n24277) );
  NOR2XL U3422 ( .A(n5914), .B(n3771), .Y(n3770) );
  XNOR2X2 U3423 ( .A(n5209), .B(n5208), .Y(n23522) );
  NAND3X1 U3424 ( .A(n5453), .B(n5451), .C(n5449), .Y(n24218) );
  XOR2X2 U3425 ( .A(n3436), .B(n5018), .Y(n5017) );
  XOR2X1 U3426 ( .A(n5920), .B(n23459), .Y(n23479) );
  XOR2X1 U3427 ( .A(n10717), .B(n10716), .Y(n3325) );
  XNOR2X1 U3428 ( .A(n10712), .B(n5479), .Y(n5478) );
  CLKINVX4 U3429 ( .A(n20425), .Y(n25300) );
  BUFX12 U3430 ( .A(n10728), .Y(n3139) );
  INVX2 U3431 ( .A(n24117), .Y(n24256) );
  OAI21XL U3432 ( .A0(n4788), .A1(n9037), .B0(n9036), .Y(n24451) );
  OAI21XL U3433 ( .A0(n3391), .A1(n24275), .B0(n3390), .Y(n5913) );
  INVX1 U3434 ( .A(n4501), .Y(n24048) );
  INVX1 U3435 ( .A(n4767), .Y(n4768) );
  XOR2X1 U3436 ( .A(n4967), .B(n3737), .Y(n24160) );
  NOR2X2 U3437 ( .A(n24031), .B(n24030), .Y(n25778) );
  XOR2X1 U3438 ( .A(n4296), .B(n20982), .Y(n23568) );
  NAND2X1 U3439 ( .A(n4524), .B(n3437), .Y(n3436) );
  XOR2XL U3440 ( .A(n23591), .B(n23590), .Y(n23626) );
  XOR2X1 U3441 ( .A(n20896), .B(n20895), .Y(n20908) );
  XOR2X1 U3442 ( .A(n20281), .B(n20280), .Y(n23612) );
  XOR2X1 U3443 ( .A(n20859), .B(n20858), .Y(n3483) );
  XOR2X1 U3444 ( .A(n23538), .B(n23537), .Y(n23611) );
  OAI2BB1X1 U3445 ( .A0N(n5969), .A1N(n21045), .B0(n5968), .Y(n3976) );
  XOR2X1 U3446 ( .A(n20332), .B(n20331), .Y(n4155) );
  XOR2X1 U3447 ( .A(n5254), .B(n23496), .Y(n23926) );
  XOR2X1 U3448 ( .A(n20971), .B(n21030), .Y(n5312) );
  XOR2X1 U3449 ( .A(n20285), .B(n20616), .Y(n20620) );
  OAI21X2 U3450 ( .A0(n4059), .A1(n23748), .B0(n4058), .Y(n23751) );
  NOR2X1 U3451 ( .A(n5030), .B(n3140), .Y(n5900) );
  NAND2X2 U3452 ( .A(n3137), .B(n25796), .Y(n3646) );
  XOR2X1 U3453 ( .A(n21021), .B(n21020), .Y(n24135) );
  XOR2X1 U3454 ( .A(n4293), .B(n4292), .Y(n23569) );
  XOR2X1 U3455 ( .A(n20758), .B(n20815), .Y(n20819) );
  XOR2X1 U3456 ( .A(n20871), .B(n20870), .Y(n20900) );
  NOR2X1 U3457 ( .A(n5353), .B(n5352), .Y(n5351) );
  XOR2X1 U3458 ( .A(n3877), .B(n4122), .Y(n4000) );
  NAND3BXL U3459 ( .AN(n23565), .B(n5429), .C(n3015), .Y(n3409) );
  NOR2X1 U3460 ( .A(n25127), .B(n4174), .Y(n4173) );
  BUFX3 U3461 ( .A(n25201), .Y(n22486) );
  CLKINVX3 U3462 ( .A(n20194), .Y(n24908) );
  BUFX12 U3463 ( .A(n5211), .Y(n4267) );
  CLKINVX2 U3464 ( .A(n4621), .Y(n4788) );
  CLKINVX4 U3465 ( .A(n19043), .Y(n4215) );
  CLKINVX3 U3466 ( .A(n5914), .Y(n5911) );
  INVX1 U3467 ( .A(n15935), .Y(n24775) );
  NOR2X1 U3468 ( .A(n3014), .B(n5033), .Y(n5429) );
  INVX1 U3469 ( .A(n19103), .Y(n5191) );
  XOR2X1 U3470 ( .A(n5483), .B(n3142), .Y(n23723) );
  OAI21X2 U3471 ( .A0(n23748), .A1(n5977), .B0(n13037), .Y(n4058) );
  NAND2X2 U3472 ( .A(n3657), .B(n3971), .Y(n4501) );
  NAND2X1 U3473 ( .A(n14643), .B(n3083), .Y(n23743) );
  XNOR2X1 U3474 ( .A(n23744), .B(n20676), .Y(n23592) );
  NOR2X1 U3475 ( .A(n4053), .B(n4052), .Y(n4063) );
  NAND2X1 U3476 ( .A(n4061), .B(n4060), .Y(n4059) );
  NAND3X1 U3477 ( .A(n4218), .B(n4217), .C(n4216), .Y(n24178) );
  XNOR2X1 U3478 ( .A(n23734), .B(n4395), .Y(n24057) );
  NOR2BX1 U3479 ( .AN(n3627), .B(n23635), .Y(n5062) );
  INVX1 U3480 ( .A(n19019), .Y(n19050) );
  INVX1 U3481 ( .A(n3132), .Y(n3078) );
  NAND3X2 U3482 ( .A(n5978), .B(n3760), .C(n3759), .Y(n23748) );
  NAND2BX2 U3483 ( .AN(n4093), .B(n4094), .Y(n5917) );
  INVX4 U3484 ( .A(n6106), .Y(n3137) );
  NAND2BX1 U3485 ( .AN(n3627), .B(n23641), .Y(n5700) );
  AOI21X1 U3486 ( .A0(n24064), .A1(n24063), .B0(n3215), .Y(n24071) );
  INVX1 U3487 ( .A(n5364), .Y(n7871) );
  NOR2X1 U3488 ( .A(n20756), .B(n20760), .Y(n3596) );
  NOR2X1 U3489 ( .A(n4867), .B(n24041), .Y(n3971) );
  BUFX8 U3490 ( .A(n23738), .Y(n3132) );
  INVX1 U3491 ( .A(n20697), .Y(n3015) );
  INVX2 U3492 ( .A(n23709), .Y(n3083) );
  NAND2BX2 U3493 ( .AN(n17427), .B(n3849), .Y(n24262) );
  NOR2X2 U3494 ( .A(n4855), .B(n17425), .Y(n17433) );
  INVXL U3495 ( .A(n3351), .Y(n3337) );
  INVX1 U3496 ( .A(n17464), .Y(n20923) );
  NOR2X1 U3497 ( .A(n8996), .B(n8995), .Y(n20384) );
  NAND2X1 U3498 ( .A(n5438), .B(n3837), .Y(n4093) );
  NOR2X1 U3499 ( .A(n5698), .B(n3329), .Y(n3336) );
  NOR2X1 U3500 ( .A(n5848), .B(n17394), .Y(n4142) );
  NAND2X1 U3501 ( .A(n3851), .B(n4105), .Y(n20693) );
  AND2X2 U3502 ( .A(n17413), .B(n24259), .Y(n3849) );
  INVX2 U3503 ( .A(n17423), .Y(n17432) );
  AND2X1 U3504 ( .A(n4198), .B(n5439), .Y(n4244) );
  INVX1 U3505 ( .A(n5834), .Y(n4855) );
  INVX1 U3506 ( .A(n5989), .Y(n4867) );
  INVX1 U3507 ( .A(n5500), .Y(n4474) );
  INVX1 U3508 ( .A(n4994), .Y(n13038) );
  INVX1 U3509 ( .A(n17463), .Y(n20931) );
  INVX1 U3510 ( .A(n20926), .Y(n5750) );
  INVXL U3511 ( .A(n4597), .Y(n3723) );
  NAND2BX2 U3512 ( .AN(n5306), .B(n3011), .Y(n20707) );
  NOR2XL U3513 ( .A(n17431), .B(n23639), .Y(n3425) );
  NAND2X2 U3514 ( .A(n4581), .B(n21110), .Y(n25542) );
  NOR2XL U3515 ( .A(n4579), .B(cs[2]), .Y(n24288) );
  INVX1 U3516 ( .A(n3852), .Y(n3851) );
  NAND2XL U3517 ( .A(n5281), .B(n5074), .Y(n4191) );
  NOR2BXL U3518 ( .AN(n5174), .B(n20638), .Y(n5173) );
  OAI2BB1X1 U3519 ( .A0N(n20402), .A1N(n9032), .B0(n9031), .Y(n20379) );
  NOR2X1 U3520 ( .A(n5933), .B(n24044), .Y(n5932) );
  NOR2X1 U3521 ( .A(n4198), .B(n19023), .Y(n4023) );
  OAI21X1 U3522 ( .A0(n23957), .A1(n15784), .B0(n15783), .Y(n23959) );
  AND2X2 U3523 ( .A(n5989), .B(n4656), .Y(n4597) );
  CLKINVX3 U3524 ( .A(n17482), .Y(n23739) );
  INVX2 U3525 ( .A(n3450), .Y(n4476) );
  NAND2X2 U3526 ( .A(n3545), .B(n20865), .Y(n20760) );
  AOI2BB2X1 U3527 ( .B0(n20121), .B1(n20120), .A0N(n20120), .A1N(n20121), .Y(
        n24389) );
  NOR2X2 U3528 ( .A(n3604), .B(n5602), .Y(n19059) );
  NAND2X1 U3529 ( .A(n17463), .B(n17467), .Y(n17359) );
  NAND2X2 U3530 ( .A(n5216), .B(n20642), .Y(n5074) );
  AOI21X2 U3531 ( .A0(n5741), .A1(n10718), .B0(n5740), .Y(n19053) );
  AOI21X1 U3532 ( .A0(n4159), .A1(n5499), .B0(n14663), .Y(n20677) );
  NOR2X2 U3533 ( .A(n23733), .B(n3147), .Y(n5446) );
  NOR2X2 U3534 ( .A(n21037), .B(n3144), .Y(n3910) );
  NAND2BX1 U3535 ( .AN(n23634), .B(n17203), .Y(n23641) );
  OAI21XL U3536 ( .A0(n14724), .A1(n24034), .B0(n24029), .Y(n5500) );
  NAND2XL U3537 ( .A(n15786), .B(n15781), .Y(n23957) );
  NOR2XL U3538 ( .A(n20380), .B(n9026), .Y(n9032) );
  NOR2X1 U3539 ( .A(n23433), .B(n23442), .Y(n19090) );
  NOR2X1 U3540 ( .A(n20663), .B(n23711), .Y(n5389) );
  NOR2X1 U3541 ( .A(n20170), .B(n20166), .Y(n24064) );
  BUFX3 U3542 ( .A(n10736), .Y(n10727) );
  INVX1 U3543 ( .A(n14661), .Y(n23442) );
  NAND2X2 U3544 ( .A(n4306), .B(n17482), .Y(n3318) );
  NAND2X1 U3545 ( .A(n23485), .B(n23484), .Y(n23486) );
  INVX1 U3546 ( .A(n14668), .Y(n23433) );
  INVX1 U3547 ( .A(n14688), .Y(n23711) );
  NAND3X1 U3548 ( .A(n5437), .B(n18973), .C(n5919), .Y(n4374) );
  NOR2X2 U3549 ( .A(n3871), .B(n4986), .Y(n23436) );
  NAND2BX2 U3550 ( .AN(n18977), .B(n18978), .Y(n3444) );
  INVX1 U3551 ( .A(n14724), .Y(n3143) );
  NAND3X1 U3552 ( .A(n5499), .B(n4159), .C(n14663), .Y(n20678) );
  NOR2X1 U3553 ( .A(n5318), .B(n3142), .Y(n5317) );
  AOI2BB1X1 U3554 ( .A0N(n25138), .A1N(n15770), .B0(n15769), .Y(n15786) );
  XNOR2X1 U3555 ( .A(n17369), .B(n17368), .Y(n17470) );
  AOI2BB1X2 U3556 ( .A0N(n23272), .A1N(n22200), .B0(n22199), .Y(n22217) );
  XNOR2X2 U3557 ( .A(n3932), .B(n4598), .Y(n17466) );
  OAI21XL U3558 ( .A0(n25301), .A1(n9014), .B0(n9013), .Y(n20380) );
  OAI21XL U3559 ( .A0(n24462), .A1(n20155), .B0(n20154), .Y(n20170) );
  AND2X2 U3560 ( .A(n23495), .B(n10703), .Y(n4648) );
  OAI21XL U3561 ( .A0(n19014), .A1(n18995), .B0(n18994), .Y(n18998) );
  CLKINVX3 U3562 ( .A(n5499), .Y(n14724) );
  XOR2X1 U3563 ( .A(n5237), .B(n10178), .Y(n17483) );
  INVX1 U3564 ( .A(n19099), .Y(n17481) );
  INVX1 U3565 ( .A(n4077), .Y(n4076) );
  NAND3BX2 U3566 ( .AN(n7319), .B(n20618), .C(n20762), .Y(n3520) );
  OAI2BB1X1 U3567 ( .A0N(n17353), .A1N(n3781), .B0(n5054), .Y(n5660) );
  NAND2XL U3568 ( .A(n20277), .B(n20278), .Y(n3534) );
  OAI21X2 U3569 ( .A0(n17382), .A1(n3335), .B0(n5058), .Y(n4161) );
  XOR2X1 U3570 ( .A(n19018), .B(n4697), .Y(n20701) );
  NOR2X1 U3571 ( .A(n4983), .B(n4982), .Y(n4416) );
  OAI2BB1XL U3572 ( .A0N(n10710), .A1N(n10709), .B0(n20944), .Y(n10711) );
  NOR2BXL U3573 ( .AN(n17452), .B(n17235), .Y(n3933) );
  NOR2X1 U3574 ( .A(n24804), .B(n23200), .Y(n24462) );
  NOR2X1 U3575 ( .A(n20538), .B(n8997), .Y(n25301) );
  NOR2X1 U3576 ( .A(n18830), .B(n6030), .Y(n5919) );
  AOI21X1 U3577 ( .A0(n5498), .A1(n5497), .B0(n4160), .Y(n4159) );
  OAI21XL U3578 ( .A0(n17365), .A1(n3335), .B0(n17364), .Y(n17369) );
  XOR2X2 U3579 ( .A(n10602), .B(n4687), .Y(n20273) );
  XOR2X2 U3580 ( .A(n4368), .B(n12850), .Y(n20312) );
  XOR2X2 U3581 ( .A(n3470), .B(n4615), .Y(n13028) );
  XOR2X2 U3582 ( .A(n4202), .B(n18856), .Y(n19020) );
  XOR2X2 U3583 ( .A(n5890), .B(n4596), .Y(n19044) );
  XOR2X2 U3584 ( .A(n3430), .B(n18860), .Y(n18978) );
  XOR2X2 U3585 ( .A(n12813), .B(n4686), .Y(n13025) );
  XOR2X2 U3586 ( .A(n6110), .B(n4695), .Y(n4994) );
  XNOR2X2 U3587 ( .A(n17340), .B(n4632), .Y(n17435) );
  XOR2X2 U3588 ( .A(n3311), .B(n4625), .Y(n17480) );
  XOR2X2 U3589 ( .A(n4859), .B(n4628), .Y(n4306) );
  XOR2X2 U3590 ( .A(n4516), .B(n12806), .Y(n23749) );
  CLKINVX3 U3591 ( .A(n15638), .Y(n3076) );
  INVX2 U3592 ( .A(n13029), .Y(n5410) );
  CLKINVX3 U3593 ( .A(n23460), .Y(n3033) );
  OAI21XL U3594 ( .A0(n17305), .A1(n17251), .B0(n17250), .Y(n17256) );
  CLKINVX3 U3595 ( .A(n6058), .Y(n4442) );
  NAND4X1 U3596 ( .A(n20665), .B(n14687), .C(n14686), .D(n14685), .Y(n14691)
         );
  NAND2X1 U3597 ( .A(n23588), .B(n23589), .Y(n20983) );
  NOR2BX2 U3598 ( .AN(n12797), .B(n4517), .Y(n4516) );
  OAI21X2 U3599 ( .A0(n12811), .A1(n3415), .B0(n4050), .Y(n12813) );
  INVX1 U3600 ( .A(n17356), .Y(n5054) );
  OAI21X2 U3601 ( .A0(n3415), .A1(n12834), .B0(n12851), .Y(n3470) );
  NAND2X1 U3602 ( .A(n7834), .B(n7833), .Y(n7835) );
  NAND2X1 U3603 ( .A(n20330), .B(n20327), .Y(n20972) );
  OAI21X2 U3604 ( .A0(n19014), .A1(n18861), .B0(n18862), .Y(n3430) );
  OAI21X1 U3605 ( .A0(n5237), .A1(n10446), .B0(n10464), .Y(n10322) );
  OAI21X2 U3606 ( .A0(n3415), .A1(n12828), .B0(n4493), .Y(n4379) );
  OAI21X2 U3607 ( .A0(n3415), .A1(n12861), .B0(n12860), .Y(n3884) );
  OAI21X2 U3608 ( .A0(n19014), .A1(n18950), .B0(n18949), .Y(n3399) );
  NAND2X1 U3609 ( .A(n3334), .B(n17336), .Y(n17340) );
  OAI21X1 U3610 ( .A0(n5237), .A1(n10629), .B0(n10628), .Y(n10633) );
  NAND3BXL U3611 ( .AN(n14662), .B(n23447), .C(n20980), .Y(n14666) );
  AOI21X2 U3612 ( .A0(n6175), .A1(n3948), .B0(n3947), .Y(n17413) );
  XOR2X1 U3613 ( .A(n7813), .B(n4691), .Y(n20282) );
  XOR2X1 U3614 ( .A(n10216), .B(n4602), .Y(n20988) );
  XOR2X1 U3615 ( .A(n10225), .B(n4605), .Y(n4331) );
  XOR2X1 U3616 ( .A(n4812), .B(n4589), .Y(n19048) );
  OAI2BB1X1 U3617 ( .A0N(n5249), .A1N(n5248), .B0(n3274), .Y(n3273) );
  XNOR2X1 U3618 ( .A(n3949), .B(n17248), .Y(n17445) );
  OAI21X1 U3619 ( .A0(n19014), .A1(n19013), .B0(n19012), .Y(n19018) );
  XNOR2X1 U3620 ( .A(n14508), .B(n14507), .Y(n14684) );
  AOI21X1 U3621 ( .A0(n3781), .A1(n4943), .B0(n4942), .Y(n3795) );
  XNOR2X1 U3622 ( .A(n7700), .B(n7699), .Y(n20363) );
  XNOR2X1 U3623 ( .A(n7804), .B(n7803), .Y(n20369) );
  XNOR2X1 U3624 ( .A(n14572), .B(n14571), .Y(n14668) );
  XNOR2X1 U3625 ( .A(n14492), .B(n14491), .Y(n23706) );
  OAI21X1 U3626 ( .A0(n5237), .A1(n10484), .B0(n10483), .Y(n3309) );
  XOR2X2 U3627 ( .A(n3551), .B(n4610), .Y(n20816) );
  XOR2X2 U3628 ( .A(n4366), .B(n12857), .Y(n13026) );
  XOR2X1 U3629 ( .A(n4071), .B(n10611), .Y(n19099) );
  XOR2X1 U3630 ( .A(n3394), .B(n17228), .Y(n17455) );
  OAI21XL U3631 ( .A0(n10243), .A1(n10179), .B0(n10182), .Y(n10225) );
  OAI21XL U3632 ( .A0(n3494), .A1(n7795), .B0(n7794), .Y(n7804) );
  OAI21XL U3633 ( .A0(n10243), .A1(n10218), .B0(n10217), .Y(n10222) );
  OAI21XL U3634 ( .A0(n17305), .A1(n17244), .B0(n17243), .Y(n3949) );
  OAI21XL U3635 ( .A0(n14677), .A1(n14676), .B0(n14675), .Y(n14681) );
  OAI21XL U3636 ( .A0(n14677), .A1(n14505), .B0(n14504), .Y(n14508) );
  OAI21XL U3637 ( .A0(n10656), .A1(n10606), .B0(n10605), .Y(n4812) );
  OAI21XL U3638 ( .A0(n10236), .A1(n10243), .B0(n10235), .Y(n5139) );
  OAI21XL U3639 ( .A0(n18869), .A1(n18925), .B0(n18868), .Y(n18872) );
  INVXL U3640 ( .A(n17265), .Y(n3948) );
  OAI21XL U3641 ( .A0(n10243), .A1(n10212), .B0(n10211), .Y(n10216) );
  OAI21XL U3642 ( .A0(n14677), .A1(n14554), .B0(n14553), .Y(n14558) );
  INVX1 U3643 ( .A(n10642), .Y(n10483) );
  INVX1 U3644 ( .A(n10738), .Y(n19077) );
  INVX1 U3645 ( .A(n10737), .Y(n20893) );
  NOR2X2 U3646 ( .A(n3415), .B(n12798), .Y(n4517) );
  OR2X2 U3647 ( .A(n4917), .B(n3469), .Y(n4378) );
  OAI21X2 U3648 ( .A0(n5237), .A1(n10655), .B0(n10654), .Y(n5474) );
  XOR2X1 U3649 ( .A(n3494), .B(n7307), .Y(n20853) );
  OAI21X2 U3650 ( .A0(n3415), .A1(n12855), .B0(n12854), .Y(n4366) );
  NOR2X2 U3651 ( .A(n24259), .B(n17294), .Y(n3947) );
  XOR2X1 U3652 ( .A(n4405), .B(n18908), .Y(n23456) );
  XOR2X1 U3653 ( .A(n12929), .B(n12878), .Y(n20317) );
  XOR2X1 U3654 ( .A(n10246), .B(n4603), .Y(n6058) );
  XOR2X1 U3655 ( .A(n4011), .B(n12932), .Y(n21017) );
  OAI21X1 U3656 ( .A0(n14677), .A1(n14513), .B0(n14512), .Y(n14518) );
  XOR2X1 U3657 ( .A(n3885), .B(n12900), .Y(n20315) );
  XNOR2X1 U3658 ( .A(n7486), .B(n7485), .Y(n20869) );
  AOI21X1 U3659 ( .A0(n12865), .A1(n12827), .B0(n12826), .Y(n4493) );
  OAI21XL U3660 ( .A0(n14677), .A1(n14489), .B0(n14488), .Y(n14492) );
  XNOR2X1 U3661 ( .A(n14501), .B(n14500), .Y(n14688) );
  OAI21X1 U3662 ( .A0(n17305), .A1(n17225), .B0(n17226), .Y(n3394) );
  XOR2X2 U3663 ( .A(n3881), .B(n12877), .Y(n13036) );
  AOI21X1 U3664 ( .A0(n12974), .A1(n12977), .B0(n12868), .Y(n4123) );
  OAI21XL U3665 ( .A0(n14677), .A1(n14498), .B0(n14497), .Y(n14501) );
  OAI21XL U3666 ( .A0(n14677), .A1(n14562), .B0(n14561), .Y(n14566) );
  OAI21XL U3667 ( .A0(n14638), .A1(n14617), .B0(n14616), .Y(n14622) );
  OAI21XL U3668 ( .A0(n10619), .A1(n10618), .B0(n10617), .Y(n10627) );
  INVX4 U3669 ( .A(n20066), .Y(n3075) );
  CLKINVX4 U3670 ( .A(n15688), .Y(n3077) );
  OAI21XL U3671 ( .A0(n18925), .A1(n18906), .B0(n18905), .Y(n4405) );
  OAI21XL U3672 ( .A0(n14638), .A1(n14631), .B0(n14630), .Y(n14635) );
  INVX1 U3673 ( .A(n18717), .Y(n18718) );
  OAI21X2 U3674 ( .A0(n3708), .A1(n3422), .B0(n17213), .Y(n5091) );
  NOR2X1 U3675 ( .A(n4411), .B(n4433), .Y(n3345) );
  NAND2BX2 U3676 ( .AN(n4003), .B(n3985), .Y(n3843) );
  AOI2BB1X1 U3677 ( .A0N(n17204), .A1N(n17257), .B0(n17259), .Y(n17264) );
  OAI2BB1X1 U3678 ( .A0N(n18829), .A1N(n6182), .B0(n6029), .Y(n18830) );
  NAND2BX1 U3679 ( .AN(n18716), .B(n19007), .Y(n18719) );
  OAI21X1 U3680 ( .A0(n14533), .A1(n14350), .B0(n5493), .Y(n14351) );
  XOR2X1 U3681 ( .A(n3587), .B(n7318), .Y(n10739) );
  OAI2BB1XL U3682 ( .A0N(n10281), .A1N(n10282), .B0(n10280), .Y(n4329) );
  OAI21X1 U3683 ( .A0(n14677), .A1(n14524), .B0(n14523), .Y(n14528) );
  OAI22X2 U3684 ( .A0(n3713), .A1(n12972), .B0(n23484), .B1(n12971), .Y(n3748)
         );
  NOR2BX2 U3685 ( .AN(n8936), .B(n8934), .Y(n8997) );
  NAND2XL U3686 ( .A(n12992), .B(n4700), .Y(n3984) );
  OAI21X1 U3687 ( .A0(n3380), .A1(n12879), .B0(n3649), .Y(n3881) );
  XNOR2X1 U3688 ( .A(n7451), .B(n7450), .Y(n20277) );
  OAI21XL U3689 ( .A0(n12929), .A1(n12885), .B0(n12884), .Y(n4021) );
  XOR2X2 U3690 ( .A(n3708), .B(n17215), .Y(n24259) );
  XOR2X2 U3691 ( .A(n4327), .B(n10207), .Y(n20944) );
  XOR2X2 U3692 ( .A(n4481), .B(n13648), .Y(n23481) );
  XNOR2X2 U3693 ( .A(n17305), .B(n17212), .Y(n20692) );
  XOR2X2 U3694 ( .A(n18925), .B(n18924), .Y(n6024) );
  XOR2X1 U3695 ( .A(n4543), .B(n7441), .Y(n20278) );
  CLKINVX3 U3696 ( .A(n3129), .Y(n22426) );
  CLKINVX3 U3697 ( .A(n14476), .Y(n14638) );
  OAI21XL U3698 ( .A0(n7446), .A1(n7423), .B0(n7445), .Y(n3587) );
  AND2X1 U3699 ( .A(n13647), .B(n13980), .Y(n13648) );
  OAI21XL U3700 ( .A0(n18984), .A1(n18716), .B0(n18715), .Y(n18717) );
  INVXL U3701 ( .A(n12865), .Y(n4080) );
  INVX1 U3702 ( .A(n12974), .Y(n4079) );
  OAI21XL U3703 ( .A0(n3126), .A1(n23223), .B0(n22187), .Y(n22192) );
  NAND2X1 U3704 ( .A(n4351), .B(n4350), .Y(n6070) );
  OAI2BB1X1 U3705 ( .A0N(n7437), .A1N(n7311), .B0(n7310), .Y(n7316) );
  BUFX3 U3706 ( .A(n9003), .Y(n20597) );
  NAND2X1 U3707 ( .A(n3567), .B(n7322), .Y(n3566) );
  NAND2BXL U3708 ( .AN(n7421), .B(n3569), .Y(n3568) );
  OAI21XL U3709 ( .A0(n12891), .A1(n12906), .B0(n12907), .Y(n4433) );
  AOI21X1 U3710 ( .A0(n14672), .A1(n14679), .B0(n14349), .Y(n5493) );
  INVX1 U3711 ( .A(n24917), .Y(n15745) );
  OAI21XL U3712 ( .A0(n14567), .A1(n14521), .B0(n14520), .Y(n14560) );
  CLKINVX4 U3713 ( .A(n22343), .Y(n3129) );
  INVX1 U3714 ( .A(n24250), .Y(n6030) );
  NAND2X1 U3715 ( .A(n3649), .B(n12880), .Y(n12881) );
  NOR2X1 U3716 ( .A(n20078), .B(n19897), .Y(n20065) );
  NOR2X1 U3717 ( .A(n15700), .B(n15517), .Y(n15687) );
  INVX1 U3718 ( .A(n19007), .Y(n4248) );
  NAND2X1 U3719 ( .A(n13000), .B(n12999), .Y(n4700) );
  NOR2X1 U3720 ( .A(n22136), .B(n21957), .Y(n22123) );
  NAND2X1 U3721 ( .A(n12990), .B(n4313), .Y(n12992) );
  NAND2X1 U3722 ( .A(n4055), .B(n12867), .Y(n12974) );
  NAND2XL U3723 ( .A(n14673), .B(n14679), .Y(n14350) );
  AOI21X1 U3724 ( .A0(n17122), .A1(n17321), .B0(n17121), .Y(n17123) );
  OAI21X1 U3725 ( .A0(n14502), .A1(n14346), .B0(n14345), .Y(n14672) );
  ADDFHX1 U3726 ( .A(n18767), .B(n23638), .CI(n17184), .CO(n23637), .S(n25136)
         );
  CLKINVX3 U3727 ( .A(n3072), .Y(n3032) );
  OAI21XL U3728 ( .A0(n3067), .A1(n20445), .B0(n8998), .Y(n20392) );
  INVX1 U3729 ( .A(n10200), .Y(n3151) );
  AOI2BB2X1 U3730 ( .B0(n24042), .B1(n24043), .A0N(n24043), .A1N(n24042), .Y(
        n24040) );
  NAND2X2 U3731 ( .A(n12780), .B(n12978), .Y(n12985) );
  NOR2X2 U3732 ( .A(n4104), .B(n3328), .Y(n17124) );
  OAI21XL U3733 ( .A0(n19008), .A1(n19015), .B0(n19016), .Y(n18993) );
  INVX1 U3734 ( .A(n5638), .Y(n5338) );
  NAND2X1 U3735 ( .A(n17239), .B(n16866), .Y(n3361) );
  OAI21X2 U3736 ( .A0(n18857), .A1(n18862), .B0(n18858), .Y(n18928) );
  NAND2BX1 U3737 ( .AN(n12991), .B(n12865), .Y(n4313) );
  NOR2X1 U3738 ( .A(n8948), .B(n8768), .Y(n8936) );
  CLKINVX4 U3739 ( .A(n25273), .Y(n3127) );
  AOI2BB1X2 U3740 ( .A0N(n10604), .A1N(n10479), .B0(n4364), .Y(n4363) );
  NAND2X1 U3741 ( .A(n18677), .B(n18676), .Y(n18858) );
  NOR2X2 U3742 ( .A(n16859), .B(n16858), .Y(n17227) );
  CLKINVX3 U3743 ( .A(n15764), .Y(n25271) );
  NAND2X1 U3744 ( .A(n17107), .B(n17106), .Y(n17314) );
  INVX1 U3745 ( .A(n22250), .Y(n22395) );
  NOR2X1 U3746 ( .A(n10175), .B(n10176), .Y(n10446) );
  OAI21XL U3747 ( .A0(n3030), .A1(n20083), .B0(n20152), .Y(n20202) );
  OAI21XL U3748 ( .A0(n10556), .A1(n10637), .B0(n5256), .Y(n10576) );
  NOR2BX1 U3749 ( .AN(n17111), .B(n5055), .Y(n17327) );
  AOI21X2 U3750 ( .A0(n4408), .A1(n3761), .B0(n3367), .Y(n18400) );
  NOR2X2 U3751 ( .A(n17237), .B(n17245), .Y(n16866) );
  NOR2X2 U3752 ( .A(n12981), .B(n12980), .Y(n12978) );
  NOR2X2 U3753 ( .A(n10218), .B(n10219), .Y(n10240) );
  NOR2X2 U3754 ( .A(n17257), .B(n17260), .Y(n17206) );
  OAI21X2 U3755 ( .A0(n17220), .A1(n17253), .B0(n17221), .Y(n3362) );
  OAI21X2 U3756 ( .A0(n17299), .A1(n17295), .B0(n17300), .Y(n17239) );
  OAI21X2 U3757 ( .A0(n10464), .A1(n10465), .B0(n10463), .Y(n10503) );
  OAI21X1 U3758 ( .A0(n14545), .A1(n14541), .B0(n14546), .Y(n14534) );
  NOR2X2 U3759 ( .A(n16853), .B(n16852), .Y(n17231) );
  NAND2X1 U3760 ( .A(n10141), .B(n10140), .Y(n10230) );
  NOR2X2 U3761 ( .A(n18676), .B(n18677), .Y(n18857) );
  NAND2X2 U3762 ( .A(n16846), .B(n16847), .Y(n17213) );
  NOR2X2 U3763 ( .A(n12764), .B(n12763), .Y(n12980) );
  NAND2X1 U3764 ( .A(n16853), .B(n16852), .Y(n17232) );
  NAND2X2 U3765 ( .A(n16851), .B(n16850), .Y(n17229) );
  NAND2X2 U3766 ( .A(n10128), .B(n10129), .Y(n10217) );
  NOR2X2 U3767 ( .A(n16864), .B(n16865), .Y(n17245) );
  NAND2X2 U3768 ( .A(n18402), .B(n18401), .Y(n4507) );
  NAND2X1 U3769 ( .A(n16856), .B(n16857), .Y(n17221) );
  NAND2X2 U3770 ( .A(n16859), .B(n16858), .Y(n17295) );
  NOR2X1 U3771 ( .A(n16843), .B(n16842), .Y(n17257) );
  NOR2X2 U3772 ( .A(n16863), .B(n16862), .Y(n17237) );
  NAND2X1 U3773 ( .A(n14312), .B(n14311), .Y(n14574) );
  NAND2X1 U3774 ( .A(n18412), .B(n18413), .Y(n18891) );
  NOR2X2 U3775 ( .A(n10133), .B(n10132), .Y(n10208) );
  NAND2X1 U3776 ( .A(n18415), .B(n18414), .Y(n18875) );
  NAND2X1 U3777 ( .A(n10120), .B(n10119), .Y(n10284) );
  NOR2X2 U3778 ( .A(n10122), .B(n10121), .Y(n10200) );
  NAND2X1 U3779 ( .A(n16843), .B(n16842), .Y(n17258) );
  INVX1 U3780 ( .A(n3609), .Y(n3608) );
  NAND2BX1 U3781 ( .AN(n17112), .B(n5056), .Y(n17331) );
  NOR2BX2 U3782 ( .AN(n10466), .B(n3150), .Y(n10608) );
  NOR2X2 U3783 ( .A(n12886), .B(n12930), .Y(n12504) );
  NAND2BX1 U3784 ( .AN(n17111), .B(n5055), .Y(n17328) );
  OAI21XL U3785 ( .A0(n18703), .A1(n18956), .B0(n18702), .Y(n18981) );
  NAND2X2 U3786 ( .A(n7320), .B(n3549), .Y(n7423) );
  OAI21XL U3787 ( .A0(n5663), .A1(n5662), .B0(n5661), .Y(n17109) );
  NOR2X2 U3788 ( .A(n7317), .B(n7429), .Y(n7443) );
  NAND2X1 U3789 ( .A(n10478), .B(n4619), .Y(n10479) );
  OAI21X2 U3790 ( .A0(n12874), .A1(n3649), .B0(n12875), .Y(n3718) );
  NAND2X1 U3791 ( .A(n14629), .B(n5210), .Y(n14624) );
  NAND2XL U3792 ( .A(n7807), .B(n7812), .Y(n7681) );
  NOR2X1 U3793 ( .A(n12824), .B(n12829), .Y(n12984) );
  ADDFHX2 U3794 ( .A(n16228), .B(n16227), .CI(n16226), .CO(n16861), .S(n16859)
         );
  ADDFHX2 U3795 ( .A(n16190), .B(n16189), .CI(n16188), .CO(n16856), .S(n16855)
         );
  ADDFHX2 U3796 ( .A(n16225), .B(n16224), .CI(n16223), .CO(n16858), .S(n16857)
         );
  ADDFHX2 U3797 ( .A(n16838), .B(n16837), .CI(n16836), .CO(n16844), .S(n16843)
         );
  NAND2X2 U3798 ( .A(n12506), .B(n12505), .Y(n12907) );
  NAND2X1 U3799 ( .A(n12507), .B(n12508), .Y(n12910) );
  NAND2X1 U3800 ( .A(n7261), .B(n7260), .Y(n7313) );
  NAND2X1 U3801 ( .A(n7264), .B(n7265), .Y(n7430) );
  NOR2X1 U3802 ( .A(n18411), .B(n18410), .Y(n18886) );
  NAND2X1 U3803 ( .A(n13997), .B(n13996), .Y(n14599) );
  NOR2X2 U3804 ( .A(n10120), .B(n10119), .Y(n10283) );
  NOR2X2 U3805 ( .A(n18415), .B(n18414), .Y(n18870) );
  NAND2X1 U3806 ( .A(n13990), .B(n13989), .Y(n14619) );
  NOR2X1 U3807 ( .A(n12497), .B(n12496), .Y(n12896) );
  NOR2X1 U3808 ( .A(n18402), .B(n18401), .Y(n18923) );
  NAND2X1 U3809 ( .A(n12489), .B(n12488), .Y(n12934) );
  NAND2X1 U3810 ( .A(n18395), .B(n18394), .Y(n18732) );
  INVX1 U3811 ( .A(n17110), .Y(n5055) );
  ADDFX2 U3812 ( .A(n7852), .B(n7405), .CI(n7404), .CO(n7402), .S(n23850) );
  INVXL U3813 ( .A(n17127), .Y(n5083) );
  NOR2X1 U3814 ( .A(n7663), .B(n7664), .Y(n5396) );
  XOR2X1 U3815 ( .A(n5529), .B(n10289), .Y(n10175) );
  OAI21XL U3816 ( .A0(n12788), .A1(n12867), .B0(n5991), .Y(n12808) );
  CLKINVX3 U3817 ( .A(n9009), .Y(n3124) );
  NAND2X2 U3818 ( .A(n14526), .B(n14564), .Y(n5494) );
  NOR2X2 U3819 ( .A(n12833), .B(n4056), .Y(n12780) );
  OAI21X2 U3820 ( .A0(n3513), .A1(n6722), .B0(n3511), .Y(n3510) );
  INVX1 U3821 ( .A(n14563), .Y(n14522) );
  OAI21X2 U3822 ( .A0(n7361), .A1(n7365), .B0(n7366), .Y(n7018) );
  OAI21X2 U3823 ( .A0(n7021), .A1(n7013), .B0(n7014), .Y(n3592) );
  OAI21X2 U3824 ( .A0(n14609), .A1(n14625), .B0(n14610), .Y(n14594) );
  NOR2X2 U3825 ( .A(n3089), .B(n3088), .Y(n14551) );
  NOR2X2 U3826 ( .A(n18731), .B(n18727), .Y(n18791) );
  NOR2X1 U3827 ( .A(n10614), .B(n10623), .Y(n10478) );
  NAND2BX1 U3828 ( .AN(n12778), .B(n4037), .Y(n4036) );
  NAND2BX1 U3829 ( .AN(n3377), .B(n3711), .Y(n3716) );
  NAND2X1 U3830 ( .A(n3306), .B(n3305), .Y(n4611) );
  OAI22X2 U3831 ( .A0(n13594), .A1(n5265), .B0(n5264), .B1(n5263), .Y(n14397)
         );
  NAND2X1 U3832 ( .A(n4252), .B(n4251), .Y(n18847) );
  ADDFHX2 U3833 ( .A(n16246), .B(n16245), .CI(n16244), .CO(n16294), .S(n16226)
         );
  ADDFHX2 U3834 ( .A(n16196), .B(n16195), .CI(n16194), .CO(n16227), .S(n16223)
         );
  ADDFHX2 U3835 ( .A(n11901), .B(n11900), .CI(n11899), .CO(n12505), .S(n12503)
         );
  ADDFHX2 U3836 ( .A(n9566), .B(n9565), .CI(n9564), .CO(n10146), .S(n9558) );
  ADDFHX2 U3837 ( .A(n9529), .B(n9528), .CI(n9527), .CO(n9559), .S(n9555) );
  ADDFHX2 U3838 ( .A(n17859), .B(n17858), .CI(n17857), .CO(n18414), .S(n18412)
         );
  ADDFHX2 U3839 ( .A(n17689), .B(n17688), .CI(n17687), .CO(n18404), .S(n18402)
         );
  ADDFHX2 U3840 ( .A(n11788), .B(n11787), .CI(n11786), .CO(n12502), .S(n12501)
         );
  INVX1 U3841 ( .A(n13593), .Y(n5264) );
  OAI21XL U3842 ( .A0(n10290), .A1(n10291), .B0(n10289), .Y(n5528) );
  XOR2X1 U3843 ( .A(n16803), .B(n3421), .Y(n16806) );
  NAND2X1 U3844 ( .A(n6906), .B(n6905), .Y(n7361) );
  XOR2X1 U3845 ( .A(n5309), .B(n9413), .Y(n10061) );
  NOR2X2 U3846 ( .A(n13997), .B(n13996), .Y(n14598) );
  NAND2X1 U3847 ( .A(n13646), .B(n13645), .Y(n13980) );
  INVXL U3848 ( .A(n18679), .Y(n4252) );
  NOR2X1 U3849 ( .A(n6958), .B(n6957), .Y(n7236) );
  NOR2X2 U3850 ( .A(n13593), .B(n13592), .Y(n13594) );
  INVXL U3851 ( .A(n13592), .Y(n5263) );
  NOR2X2 U3852 ( .A(n12765), .B(n12766), .Y(n12981) );
  OAI2BB1X1 U3853 ( .A0N(n6093), .A1N(n18588), .B0(n6092), .Y(n18591) );
  XOR2X1 U3854 ( .A(n10083), .B(n5380), .Y(n4115) );
  NAND2X1 U3855 ( .A(n12766), .B(n12765), .Y(n12982) );
  ADDFX2 U3856 ( .A(n18786), .B(n11616), .CI(n11615), .CO(n11613), .S(n24285)
         );
  NAND2X1 U3857 ( .A(n13591), .B(n13590), .Y(n5265) );
  ADDFX2 U3858 ( .A(n18776), .B(n17190), .CI(n17189), .CO(n17187), .S(n25099)
         );
  OAI21X1 U3859 ( .A0(n4304), .A1(n9268), .B0(n9369), .Y(n3829) );
  OR2X2 U3860 ( .A(n14318), .B(n14317), .Y(n14564) );
  NOR2X1 U3861 ( .A(n12424), .B(n12423), .Y(n3377) );
  NOR2XL U3862 ( .A(n13591), .B(n13590), .Y(n5258) );
  OAI2BB1X1 U3863 ( .A0N(n5689), .A1N(n16302), .B0(n5688), .Y(n17015) );
  OAI2BB1X1 U3864 ( .A0N(n17647), .A1N(n17646), .B0(n6157), .Y(n18407) );
  NOR2X1 U3865 ( .A(n10473), .B(n10474), .Y(n10614) );
  NAND2X2 U3866 ( .A(n3420), .B(n5508), .Y(n3889) );
  ADDFHX1 U3867 ( .A(n16193), .B(n16192), .CI(n16191), .CO(n16228), .S(n16225)
         );
  ADDFHX1 U3868 ( .A(n12468), .B(n12467), .CI(n12466), .CO(n12490), .S(n12489)
         );
  ADDFHX1 U3869 ( .A(n16835), .B(n16834), .CI(n16833), .CO(n16825), .S(n16836)
         );
  AOI21X2 U3870 ( .A0(n3506), .A1(n6728), .B0(n6727), .Y(n3505) );
  ADDFHX1 U3871 ( .A(n10113), .B(n10112), .CI(n10111), .CO(n10119), .S(n10118)
         );
  NAND3BX1 U3872 ( .AN(n6717), .B(n6721), .C(n5616), .Y(n6722) );
  NOR2XL U3873 ( .A(n4141), .B(n4140), .Y(n3242) );
  ADDFHX1 U3874 ( .A(n18581), .B(n18580), .CI(n18579), .CO(n18675), .S(n18416)
         );
  XNOR2X1 U3875 ( .A(n22062), .B(n22061), .Y(n22448) );
  ADDFHX2 U3876 ( .A(n7254), .B(n7253), .CI(n7252), .CO(n7259), .S(n7004) );
  ADDFHX2 U3877 ( .A(n7002), .B(n7001), .CI(n7000), .CO(n7003), .S(n6958) );
  ADDFHX2 U3878 ( .A(n13907), .B(n13906), .CI(n13905), .CO(n13994), .S(n13993)
         );
  ADDFHX2 U3879 ( .A(n6901), .B(n6900), .CI(n6899), .CO(n6911), .S(n6910) );
  ADDFX2 U3880 ( .A(n10110), .B(n10109), .CI(n10108), .CO(n10100), .S(n10111)
         );
  CMPR32X1 U3881 ( .A(n7173), .B(n7172), .C(n7171), .CO(n7206), .S(n7203) );
  CMPR32X1 U3882 ( .A(n17007), .B(n17006), .C(n17005), .CO(n17009), .S(n17011)
         );
  CMPR32X1 U3883 ( .A(n16999), .B(n16998), .C(n16997), .CO(n17031), .S(n17020)
         );
  OAI21XL U3884 ( .A0(n5903), .A1(n5902), .B0(n5901), .Y(n17856) );
  INVX1 U3885 ( .A(n12427), .Y(n5508) );
  CMPR32X1 U3886 ( .A(n7640), .B(n7639), .C(n7638), .CO(n7678), .S(n7675) );
  XOR2X1 U3887 ( .A(n16787), .B(n16786), .Y(n3794) );
  ADDFX2 U3888 ( .A(n14242), .B(n14241), .CI(n14240), .CO(n14330), .S(n14327)
         );
  INVX1 U3889 ( .A(n10053), .Y(n3091) );
  ADDFX2 U3890 ( .A(n18599), .B(n18598), .CI(n18597), .CO(n18696), .S(n18687)
         );
  OAI2BB1X1 U3891 ( .A0N(n5155), .A1N(n14185), .B0(n5154), .Y(n14203) );
  NAND2BX2 U3892 ( .AN(n6726), .B(n3516), .Y(n6728) );
  NOR2X1 U3893 ( .A(n9508), .B(n9509), .Y(n4119) );
  OAI2BB1X2 U3894 ( .A0N(n17625), .A1N(n5868), .B0(n5867), .Y(n17852) );
  OAI2BB1X2 U3895 ( .A0N(n11919), .A1N(n4426), .B0(n4972), .Y(n11963) );
  NAND2X1 U3896 ( .A(n5955), .B(n5954), .Y(n16192) );
  OAI2BB1X1 U3897 ( .A0N(n10428), .A1N(n10430), .B0(n4359), .Y(n10467) );
  OR2X2 U3898 ( .A(n12767), .B(n12768), .Y(n12858) );
  OAI21XL U3899 ( .A0(n5737), .A1(n5736), .B0(n5735), .Y(n16762) );
  ADDFHX1 U3900 ( .A(n9389), .B(n9388), .CI(n9387), .CO(n9409), .S(n9417) );
  ADDFHX1 U3901 ( .A(n16483), .B(n16482), .CI(n16481), .CO(n16775), .S(n16774)
         );
  ADDFHX1 U3902 ( .A(n10098), .B(n10097), .CI(n10096), .CO(n10083), .S(n10099)
         );
  ADDFHX1 U3903 ( .A(n13549), .B(n13548), .CI(n13547), .CO(n13592), .S(n13591)
         );
  ADDFHX1 U3904 ( .A(n18391), .B(n18390), .CI(n18389), .CO(n18394), .S(n18393)
         );
  ADDFHX1 U3905 ( .A(n16566), .B(n16565), .CI(n16564), .CO(n16767), .S(n16765)
         );
  ADDFHX1 U3906 ( .A(n7493), .B(n7492), .CI(n7491), .CO(n7520), .S(n7482) );
  NAND2X1 U3907 ( .A(n6047), .B(n6046), .Y(n13992) );
  NOR2X1 U3908 ( .A(n3481), .B(n5636), .Y(n3479) );
  NOR2X1 U3909 ( .A(n12848), .B(n12841), .Y(n12779) );
  ADDFHX1 U3910 ( .A(n18577), .B(n18576), .CI(n18575), .CO(n18680), .S(n18678)
         );
  OAI21X1 U3911 ( .A0(n5623), .A1(n6717), .B0(n6716), .Y(n3512) );
  XNOR2X1 U3912 ( .A(n8829), .B(n9027), .Y(n9030) );
  ADDFHX2 U3913 ( .A(n16480), .B(n16479), .CI(n16478), .CO(n16454), .S(n16481)
         );
  ADDFHX2 U3914 ( .A(n13885), .B(n13884), .CI(n13883), .CO(n13942), .S(n13905)
         );
  ADDFHX2 U3915 ( .A(n7123), .B(n7122), .CI(n7121), .CO(n7134), .S(n7238) );
  ADDFHX2 U3916 ( .A(n16141), .B(n16140), .CI(n16139), .CO(n16170), .S(n16137)
         );
  ADDFHX2 U3917 ( .A(n6934), .B(n6933), .CI(n6932), .CO(n7001), .S(n6955) );
  ADDFHX2 U3918 ( .A(n16504), .B(n16503), .CI(n16502), .CO(n16482), .S(n16561)
         );
  ADDFHX2 U3919 ( .A(n13814), .B(n13813), .CI(n13812), .CO(n13819), .S(n13821)
         );
  ADDFHX2 U3920 ( .A(n6981), .B(n6980), .CI(n6979), .CO(n7253), .S(n7000) );
  OAI21XL U3921 ( .A0(n16828), .A1(n16829), .B0(n16827), .Y(n3774) );
  ADDFX2 U3922 ( .A(n16307), .B(n16306), .CI(n16305), .CO(n17025), .S(n16303)
         );
  CMPR32X1 U3923 ( .A(n7120), .B(n7119), .C(n7118), .CO(n7135), .S(n7239) );
  INVX1 U3924 ( .A(n13826), .Y(n3449) );
  CMPR32X1 U3925 ( .A(n16231), .B(n16230), .C(n16229), .CO(n16263), .S(n16255)
         );
  ADDFX2 U3926 ( .A(n10150), .B(n10149), .CI(n10148), .CO(n10291), .S(n10172)
         );
  CMPR32X1 U3927 ( .A(n9554), .B(n9553), .C(n9552), .CO(n9561), .S(n9524) );
  ADDFX2 U3928 ( .A(n14239), .B(n14238), .CI(n14237), .CO(n14240), .S(n14222)
         );
  CLKINVX3 U3929 ( .A(n6732), .Y(n3481) );
  CMPR32X1 U3930 ( .A(n16292), .B(n16291), .C(n16290), .CO(n16299), .S(n16261)
         );
  OAI21XL U3931 ( .A0(n3980), .A1(n3979), .B0(n3978), .Y(n12686) );
  INVXL U3932 ( .A(n16018), .Y(n3342) );
  ADDFX2 U3933 ( .A(n14271), .B(n14270), .CI(n14269), .CO(n14273), .S(n14258)
         );
  INVX1 U3934 ( .A(n16304), .Y(n5690) );
  XOR2X1 U3935 ( .A(n5615), .B(n6893), .Y(n6902) );
  CMPR32X1 U3936 ( .A(n18631), .B(n18630), .C(n18629), .CO(n18700), .S(n18697)
         );
  XOR2X1 U3937 ( .A(n5137), .B(n6953), .Y(n6956) );
  XOR2X1 U3938 ( .A(n3729), .B(n12447), .Y(n12478) );
  CMPR32X1 U3939 ( .A(n17043), .B(n17042), .C(n17041), .CO(n17063), .S(n17048)
         );
  OAI2BB1X1 U3940 ( .A0N(n3544), .A1N(n7177), .B0(n3543), .Y(n7212) );
  INVX1 U3941 ( .A(n6725), .Y(n3516) );
  OAI2BB1X1 U3942 ( .A0N(n5930), .A1N(n12681), .B0(n5929), .Y(n12684) );
  INVXL U3943 ( .A(n12769), .Y(n5961) );
  OAI2BB1X1 U3944 ( .A0N(n5723), .A1N(n16966), .B0(n5722), .Y(n16997) );
  XNOR2X1 U3945 ( .A(n12681), .B(n5931), .Y(n12672) );
  OAI21XL U3946 ( .A0(n8882), .A1(n8834), .B0(n8828), .Y(n8829) );
  OAI21XL U3947 ( .A0(n15632), .A1(n15584), .B0(n15578), .Y(n15579) );
  OAI21XL U3948 ( .A0(n15632), .A1(n15584), .B0(n15583), .Y(n15586) );
  OAI21XL U3949 ( .A0(n22070), .A1(n22022), .B0(n22016), .Y(n22017) );
  OAI21XL U3950 ( .A0(n8882), .A1(n8834), .B0(n8833), .Y(n8836) );
  OAI21XL U3951 ( .A0(n22070), .A1(n22022), .B0(n22021), .Y(n22024) );
  XNOR2X1 U3952 ( .A(n16300), .B(n5333), .Y(n5332) );
  OAI21XL U3953 ( .A0(n18305), .A1(n18304), .B0(n18303), .Y(n18309) );
  ADDFHX1 U3954 ( .A(n10104), .B(n10103), .CI(n10102), .CO(n10096), .S(n10113)
         );
  ADDFHX1 U3955 ( .A(n18568), .B(n18567), .CI(n18566), .CO(n18573), .S(n18576)
         );
  XNOR2X2 U3956 ( .A(n5172), .B(n9518), .Y(n9508) );
  ADDFHX1 U3957 ( .A(n7170), .B(n7169), .CI(n7168), .CO(n7174), .S(n7150) );
  OAI2BB1X1 U3958 ( .A0N(n3276), .A1N(n9763), .B0(n3275), .Y(n10055) );
  ADDFHX1 U3959 ( .A(n9458), .B(n9457), .CI(n9456), .CO(n9509), .S(n9484) );
  ADDFHX1 U3960 ( .A(n16557), .B(n16556), .CI(n16555), .CO(n16562), .S(n16564)
         );
  ADDFHX1 U3961 ( .A(n17800), .B(n17799), .CI(n17798), .CO(n17847), .S(n17849)
         );
  ADDFHX1 U3962 ( .A(n14178), .B(n14177), .CI(n14176), .CO(n14318), .S(n14315)
         );
  ADDFHX1 U3963 ( .A(n14175), .B(n14174), .CI(n14173), .CO(n14316), .S(n14314)
         );
  ADDFHX1 U3964 ( .A(n9767), .B(n9765), .CI(n9766), .CO(n10053), .S(n10052) );
  XNOR2X2 U3965 ( .A(n3370), .B(n3369), .Y(n16169) );
  XNOR2X1 U3966 ( .A(n8874), .B(n8873), .Y(n20404) );
  ADDFHX1 U3967 ( .A(n16750), .B(n16749), .CI(n16748), .CO(n16752), .S(n16727)
         );
  OAI21X1 U3968 ( .A0(n4127), .A1(n4128), .B0(n3801), .Y(n3800) );
  ADDFHX1 U3969 ( .A(n9829), .B(n9828), .CI(n9827), .CO(n10051), .S(n10048) );
  XNOR2X1 U3970 ( .A(n19958), .B(n3215), .Y(n20167) );
  ADDFHX2 U3971 ( .A(n13832), .B(n13831), .CI(n13830), .CO(n13906), .S(n13824)
         );
  ADDFHX2 U3972 ( .A(n12085), .B(n12084), .CI(n12083), .CO(n12470), .S(n12086)
         );
  ADDFHX2 U3973 ( .A(n17769), .B(n17768), .CI(n17767), .CO(n17805), .S(n17842)
         );
  ADDFHX2 U3974 ( .A(n9394), .B(n9395), .CI(n9393), .CO(n9418), .S(n10063) );
  CMPR32X1 U3975 ( .A(n16814), .B(n16813), .C(n16812), .CO(n16809), .S(n16835)
         );
  CMPR32X1 U3976 ( .A(n16551), .B(n16550), .C(n16549), .CO(n16502), .S(n16566)
         );
  ADDFX2 U3977 ( .A(n16744), .B(n16743), .CI(n16742), .CO(n16734), .S(n16745)
         );
  CMPR32X1 U3978 ( .A(n18510), .B(n18509), .C(n18508), .CO(n18511), .S(n18566)
         );
  CMPR32X1 U3979 ( .A(n7188), .B(n7187), .C(n7186), .CO(n7213), .S(n7177) );
  ADDFX2 U3980 ( .A(n17821), .B(n17820), .CI(n17819), .CO(n18590), .S(n17817)
         );
  INVX1 U3981 ( .A(n17627), .Y(n5870) );
  OAI21XL U3982 ( .A0(n5775), .A1(n12476), .B0(n12475), .Y(n5774) );
  CMPR32X1 U3983 ( .A(n18456), .B(n18455), .C(n18454), .CO(n18474), .S(n18457)
         );
  CMPR32X1 U3984 ( .A(n7559), .B(n7558), .C(n7557), .CO(n7577), .S(n7560) );
  CMPR32X1 U3985 ( .A(n7200), .B(n7199), .C(n7198), .CO(n7207), .S(n7171) );
  OAI2BB1X1 U3986 ( .A0N(n6984), .A1N(n6982), .B0(n4554), .Y(n7245) );
  CMPR32X1 U3987 ( .A(n16209), .B(n16208), .C(n16207), .CO(n16229), .S(n16214)
         );
  OAI21XL U3988 ( .A0(n5292), .A1(n5291), .B0(n5290), .Y(n13812) );
  ADDFX2 U3989 ( .A(n16536), .B(n16535), .CI(n16534), .CO(n16552), .S(n16735)
         );
  OAI21XL U3990 ( .A0(n4818), .A1(n4817), .B0(n4816), .Y(n9350) );
  CMPR32X1 U3991 ( .A(n16310), .B(n16309), .C(n16308), .CO(n16993), .S(n16306)
         );
  OAI21XL U3992 ( .A0(n4870), .A1(n4869), .B0(n4868), .Y(n18371) );
  ADDFX2 U3993 ( .A(n18642), .B(n18641), .CI(n18640), .CO(n18643), .S(n18630)
         );
  ADDFX2 U3994 ( .A(n18477), .B(n18476), .CI(n18475), .CO(n18599), .S(n18487)
         );
  OAI2BB1X1 U3995 ( .A0N(n18559), .A1N(n18558), .B0(n4246), .Y(n18570) );
  CMPR32X1 U3996 ( .A(n6693), .B(n6692), .C(n6691), .CO(n6712), .S(n6673) );
  CMPR32X1 U3997 ( .A(n9808), .B(n9807), .C(n9806), .CO(n10044), .S(n10043) );
  CMPR32X1 U3998 ( .A(n3114), .B(n16206), .C(n16205), .CO(n16230), .S(n16212)
         );
  OAI21XL U3999 ( .A0(n3453), .A1(n5070), .B0(n5068), .Y(n9375) );
  OAI2BB1X1 U4000 ( .A0N(n4495), .A1N(n13500), .B0(n4494), .Y(n13522) );
  ADDFX2 U4001 ( .A(n10397), .B(n10396), .CI(n10395), .CO(n10449), .S(n10407)
         );
  XOR2X1 U4002 ( .A(n5042), .B(n16158), .Y(n16186) );
  OAI2BB1X1 U4003 ( .A0N(n4371), .A1N(n17770), .B0(n4370), .Y(n17796) );
  OAI21XL U4004 ( .A0(n20011), .A1(n19963), .B0(n19957), .Y(n19958) );
  XOR2X1 U4005 ( .A(n16448), .B(n4113), .Y(n4112) );
  OAI21XL U4006 ( .A0(n20011), .A1(n19963), .B0(n19962), .Y(n19965) );
  NAND2X1 U4007 ( .A(n3816), .B(n3815), .Y(n3814) );
  OAI21XL U4008 ( .A0(n6000), .A1(n5999), .B0(n5998), .Y(n12784) );
  XNOR2X1 U4009 ( .A(n12683), .B(n12682), .Y(n5931) );
  ADDFHX1 U4010 ( .A(n6937), .B(n6936), .CI(n6935), .CO(n6981), .S(n6933) );
  XNOR2X1 U4011 ( .A(n5041), .B(n12666), .Y(n12770) );
  ADDFHX1 U4012 ( .A(n10073), .B(n10072), .CI(n10071), .CO(n10062), .S(n10097)
         );
  ADDFHX1 U4013 ( .A(n10107), .B(n10106), .CI(n10105), .CO(n10112), .S(n10115)
         );
  ADDFHX1 U4014 ( .A(n9314), .B(n9313), .CI(n9312), .CO(n9309), .S(n9415) );
  OAI22X1 U4015 ( .A0(n4514), .A1(n4515), .B0(n3901), .B1(n3900), .Y(n3899) );
  ADDFHX1 U4016 ( .A(n13486), .B(n13485), .CI(n13484), .CO(n13548), .S(n13503)
         );
  ADDFHX1 U4017 ( .A(n16157), .B(n16156), .CI(n16155), .CO(n16193), .S(n16187)
         );
  ADDFHX1 U4018 ( .A(n16716), .B(n16715), .CI(n16714), .CO(n16749), .S(n16717)
         );
  XOR2X2 U4019 ( .A(n16415), .B(n16417), .Y(n4850) );
  ADDFHX1 U4020 ( .A(n16040), .B(n16039), .CI(n16038), .CO(n16139), .S(n16045)
         );
  ADDFHX1 U4021 ( .A(n16059), .B(n16058), .CI(n16057), .CO(n16077), .S(n16085)
         );
  ADDFHX1 U4022 ( .A(n18495), .B(n18494), .CI(n18493), .CO(n18512), .S(n18568)
         );
  ADDFHX1 U4023 ( .A(n17692), .B(n17691), .CI(n17690), .CO(n17685), .S(n18334)
         );
  ADDFHX1 U4024 ( .A(n17841), .B(n17840), .CI(n17839), .CO(n18582), .S(n17814)
         );
  ADDFHX1 U4025 ( .A(n9497), .B(n9496), .CI(n9495), .CO(n9525), .S(n9521) );
  ADDFX2 U4026 ( .A(n9300), .B(n9299), .CI(n9298), .CO(n9311), .S(n9388) );
  ADDFHX1 U4027 ( .A(n9494), .B(n9493), .CI(n9492), .CO(n9526), .S(n9518) );
  ADDFX2 U4028 ( .A(n16037), .B(n16036), .CI(n16035), .CO(n16046), .S(n16082)
         );
  ADDFHX2 U4029 ( .A(n16458), .B(n16457), .CI(n16456), .CO(n16416), .S(n16483)
         );
  ADDFHX2 U4030 ( .A(n16793), .B(n16792), .CI(n16791), .CO(n16786), .S(n16822)
         );
  ADDFHX2 U4031 ( .A(n16043), .B(n16042), .CI(n16041), .CO(n16151), .S(n16044)
         );
  ADDFHX2 U4032 ( .A(n14104), .B(n14103), .CI(n14102), .CO(n14178), .S(n14168)
         );
  OAI21XL U4033 ( .A0(n6982), .A1(n6984), .B0(n6983), .Y(n4554) );
  OAI21XL U4034 ( .A0(n16120), .A1(n16119), .B0(n16118), .Y(n3816) );
  CMPR32X1 U4035 ( .A(n13521), .B(n13520), .C(n13519), .CO(n13581), .S(n13523)
         );
  OAI21XL U4036 ( .A0(n12667), .A1(n12668), .B0(n12666), .Y(n5038) );
  CMPR32X1 U4037 ( .A(n14042), .B(n14041), .C(n14040), .CO(n14163), .S(n14066)
         );
  OAI21XL U4038 ( .A0(n13753), .A1(n13752), .B0(n13751), .Y(n5290) );
  ADDFX2 U4039 ( .A(n9380), .B(n9379), .CI(n9378), .CO(n9389), .S(n9394) );
  ADDFX2 U4040 ( .A(n16163), .B(n16162), .CI(n16161), .CO(n16215), .S(n16156)
         );
  ADDFX2 U4041 ( .A(n16443), .B(n16442), .CI(n16441), .CO(n16817), .S(n16801)
         );
  ADDFX2 U4042 ( .A(n9960), .B(n9225), .CI(n9224), .CO(n9237), .S(n9298) );
  ADDFX2 U4043 ( .A(n16106), .B(n16105), .CI(n16104), .CO(n16790), .S(n16816)
         );
  CMPR32X1 U4044 ( .A(n16525), .B(n16524), .C(n16523), .CO(n16549), .S(n16553)
         );
  CMPR32X1 U4045 ( .A(n16695), .B(n16694), .C(n16693), .CO(n16741), .S(n16715)
         );
  INVX1 U4046 ( .A(n11752), .Y(n3898) );
  ADDFX2 U4047 ( .A(n18553), .B(n18552), .CI(n18551), .CO(n18563), .S(n18561)
         );
  CMPR32X1 U4048 ( .A(n18498), .B(n18497), .C(n18496), .CO(n18494), .S(n18531)
         );
  CMPR32X1 U4049 ( .A(n6076), .B(n9235), .C(n9234), .CO(n9273), .S(n9236) );
  CMPR32X1 U4050 ( .A(n16713), .B(n16712), .C(n16711), .CO(n16718), .S(n16720)
         );
  CMPR32X1 U4051 ( .A(n16324), .B(n16323), .C(n16322), .CO(n16966), .S(n16325)
         );
  OAI21XL U4052 ( .A0(n17099), .A1(n16903), .B0(n5827), .Y(n16906) );
  INVXL U4053 ( .A(n13811), .Y(n13807) );
  ADDFX2 U4054 ( .A(n18273), .B(n18272), .CI(n18271), .CO(n18299), .S(n18293)
         );
  CMPR32X1 U4055 ( .A(n17823), .B(n17824), .C(n17822), .CO(n18556), .S(n17820)
         );
  ADDFX2 U4056 ( .A(n17789), .B(n17788), .CI(n17787), .CO(n17840), .S(n17792)
         );
  OAI2BB1X1 U4057 ( .A0N(n15995), .A1N(n15994), .B0(n5801), .Y(n16017) );
  CMPR32X1 U4058 ( .A(n12725), .B(n12724), .C(n12723), .CO(n12786), .S(n12783)
         );
  ADDFX2 U4059 ( .A(n9103), .B(n10492), .CI(n10491), .CO(n10519), .S(n10499)
         );
  ADDFX2 U4060 ( .A(n16946), .B(n16945), .CI(n16944), .CO(n16932), .S(n16968)
         );
  ADDFX2 U4061 ( .A(n18498), .B(n16936), .CI(n16935), .CO(n16933), .S(n16970)
         );
  OAI2BB1X1 U4062 ( .A0N(n5195), .A1N(n9648), .B0(n5194), .Y(n10107) );
  ADDFX2 U4063 ( .A(n9548), .B(n9547), .CI(n9546), .CO(n9587), .S(n9552) );
  ADDFX2 U4064 ( .A(n9515), .B(n9514), .CI(n9513), .CO(n9531), .S(n9520) );
  OAI21X1 U4065 ( .A0(n12431), .A1(n12432), .B0(n12430), .Y(n3650) );
  CMPR32X1 U4066 ( .A(n16912), .B(n16911), .C(n16910), .CO(n16916), .S(n16898)
         );
  CMPR32X1 U4067 ( .A(n7549), .B(n7550), .C(n7548), .CO(n7559), .S(n7543) );
  ADDFX2 U4068 ( .A(n16545), .B(n16544), .CI(n16543), .CO(n16534), .S(n16742)
         );
  OAI2BB1X1 U4069 ( .A0N(n5283), .A1N(n9823), .B0(n5282), .Y(n9807) );
  XOR2X1 U4070 ( .A(n9376), .B(n3268), .Y(n9395) );
  ADDFX2 U4071 ( .A(n16495), .B(n16494), .CI(n16493), .CO(n16490), .S(n16509)
         );
  ADDFX2 U4072 ( .A(n16896), .B(n16895), .CI(n16894), .CO(n16897), .S(n16929)
         );
  ADDFX2 U4073 ( .A(n16252), .B(n16251), .CI(n16250), .CO(n16268), .S(n16257)
         );
  OAI2BB1X1 U4074 ( .A0N(n16000), .A1N(n5808), .B0(n5807), .Y(n16036) );
  OAI2BB1X1 U4075 ( .A0N(n16090), .A1N(n3694), .B0(n3693), .Y(n16075) );
  OAI2BB1X1 U4076 ( .A0N(n11715), .A1N(n3645), .B0(n3644), .Y(n11785) );
  OAI2BB1X1 U4077 ( .A0N(n4337), .A1N(n17702), .B0(n4336), .Y(n17690) );
  XOR2X1 U4078 ( .A(n16053), .B(n3634), .Y(n16074) );
  ADDFX2 U4079 ( .A(n9467), .B(n9466), .CI(n9465), .CO(n9493), .S(n9473) );
  OAI21XL U4080 ( .A0(n4905), .A1(n4904), .B0(n4903), .Y(n12687) );
  OAI2BB1X1 U4081 ( .A0N(n9245), .A1N(n4308), .B0(n4307), .Y(n9291) );
  OAI2BB1X1 U4082 ( .A0N(n6127), .A1N(n18075), .B0(n6126), .Y(n18301) );
  OAI21XL U4083 ( .A0(n4880), .A1(n4879), .B0(n4878), .Y(n12415) );
  OAI21XL U4084 ( .A0(n4262), .A1(n4261), .B0(n4260), .Y(n13340) );
  OAI21XL U4085 ( .A0(n21970), .A1(n21969), .B0(n21968), .Y(n21971) );
  ADDFHX1 U4086 ( .A(n13489), .B(n13488), .CI(n13487), .CO(n13524), .S(n13485)
         );
  ADDFHX1 U4087 ( .A(n12063), .B(n12062), .CI(n12061), .CO(n12460), .S(n12088)
         );
  ADDFHX1 U4088 ( .A(n12456), .B(n12455), .CI(n12454), .CO(n12457), .S(n12461)
         );
  ADDFHX1 U4089 ( .A(n13627), .B(n13626), .CI(n13625), .CO(n13806), .S(n13644)
         );
  ADDFHX1 U4090 ( .A(n18098), .B(n18097), .CI(n18096), .CO(n18313), .S(n18307)
         );
  ADDFHX1 U4091 ( .A(n12042), .B(n12041), .CI(n12040), .CO(n12462), .S(n12084)
         );
  ADDFX2 U4092 ( .A(n6767), .B(n6766), .CI(n6765), .CO(n6887), .S(n6808) );
  ADDFHX1 U4093 ( .A(n13707), .B(n13706), .CI(n13705), .CO(n13743), .S(n13804)
         );
  ADDFHX1 U4094 ( .A(n11714), .B(n11713), .CI(n11712), .CO(n11769), .S(n11719)
         );
  ADDFHX1 U4095 ( .A(n16369), .B(n16368), .CI(n16367), .CO(n16434), .S(n16415)
         );
  ADDFHX1 U4096 ( .A(n12552), .B(n12551), .CI(n12550), .CO(n12566), .S(n12608)
         );
  ADDFHX1 U4097 ( .A(n10375), .B(n10374), .CI(n10373), .CO(n10394), .S(n10376)
         );
  CMPR32X1 U4098 ( .A(n12453), .B(n12452), .C(n12451), .CO(n12458), .S(n12439)
         );
  CMPR32X1 U4099 ( .A(n13937), .B(n13936), .C(n13935), .CO(n13947), .S(n13909)
         );
  CMPR32X1 U4100 ( .A(n18528), .B(n18527), .C(n18526), .CO(n18560), .S(n18583)
         );
  ADDFHX1 U4101 ( .A(n11807), .B(n11806), .CI(n11805), .CO(n11802), .S(n12476)
         );
  ADDFHX1 U4102 ( .A(n7072), .B(n7071), .CI(n7070), .CO(n7128), .S(n7125) );
  ADDFHX2 U4103 ( .A(n18343), .B(n18342), .CI(n18341), .CO(n18336), .S(n18372)
         );
  ADDFHX2 U4104 ( .A(n12438), .B(n12437), .CI(n12436), .CO(n12431), .S(n12464)
         );
  OAI21XL U4105 ( .A0(n15994), .A1(n15995), .B0(n15993), .Y(n5801) );
  ADDFX2 U4106 ( .A(n13322), .B(n13321), .CI(n13320), .CO(n13418), .S(n13336)
         );
  OAI21XL U4107 ( .A0(n12679), .A1(n12680), .B0(n12678), .Y(n4903) );
  OAI21XL U4108 ( .A0(n17609), .A1(n3169), .B0(n17608), .Y(n5477) );
  ADDFX2 U4109 ( .A(n14074), .B(n14073), .CI(n14072), .CO(n14103), .S(n14165)
         );
  ADDFX2 U4110 ( .A(n9770), .B(n9769), .CI(n9768), .CO(n9759), .S(n9831) );
  CMPR32X1 U4111 ( .A(n18074), .B(n18073), .C(n18072), .CO(n18100), .S(n18075)
         );
  CMPR32X1 U4112 ( .A(n12735), .B(n12734), .C(n12733), .CO(n12737), .S(n12724)
         );
  CMPR32X1 U4113 ( .A(n16440), .B(n16439), .C(n16438), .CO(n16802), .S(n16435)
         );
  CMPR32X1 U4114 ( .A(n12045), .B(n12044), .C(n12043), .CO(n12456), .S(n12040)
         );
  ADDFX2 U4115 ( .A(n12721), .B(n12720), .CI(n12719), .CO(n12723), .S(n12706)
         );
  CMPR32X1 U4116 ( .A(n12091), .B(n12090), .C(n12089), .CO(n12083), .S(n12113)
         );
  CMPR32X1 U4117 ( .A(n9792), .B(n9791), .C(n9790), .CO(n9787), .S(n9808) );
  CMPR32X1 U4118 ( .A(n12372), .B(n12371), .C(n12370), .CO(n12379), .S(n12378)
         );
  CMPR32X1 U4119 ( .A(n9260), .B(n9259), .C(n9258), .CO(n9285), .S(n9312) );
  CMPR32X1 U4120 ( .A(n16123), .B(n16122), .C(n16121), .CO(n16157), .S(n16118)
         );
  CMPR32X1 U4121 ( .A(n12054), .B(n12053), .C(n12052), .CO(n12441), .S(n12063)
         );
  CMPR32X1 U4122 ( .A(n16965), .B(n18525), .C(n18524), .CO(n18551), .S(n18527)
         );
  OAI21XL U4123 ( .A0(n3653), .A1(n3654), .B0(n3652), .Y(n11807) );
  OAI21XL U4124 ( .A0(n4570), .A1(n6139), .B0(n6138), .Y(n9500) );
  ADDFX2 U4125 ( .A(n11961), .B(n11960), .CI(n11959), .CO(n11968), .S(n11934)
         );
  CMPR32X1 U4126 ( .A(n10391), .B(n10390), .C(n10389), .CO(n10395), .S(n10374)
         );
  CMPR32X1 U4127 ( .A(n7233), .B(n7234), .C(n7235), .CO(n7301), .S(n7228) );
  OAI21XL U4128 ( .A0(n3287), .A1(n9435), .B0(n3303), .Y(n10076) );
  OAI21XL U4129 ( .A0(n18111), .A1(n4205), .B0(n4204), .Y(n17757) );
  ADDFX2 U4130 ( .A(n7056), .B(n6993), .CI(n6861), .CO(n7070), .S(n6961) );
  OAI21XL U4131 ( .A0(n16469), .A1(n16704), .B0(n5845), .Y(n16489) );
  ADDFX2 U4132 ( .A(n11711), .B(n11710), .CI(n11709), .CO(n11720), .S(n11789)
         );
  CMPR32X1 U4133 ( .A(n7064), .B(n7063), .C(n7062), .CO(n7106), .S(n7083) );
  ADDFX2 U4134 ( .A(n16392), .B(n16391), .CI(n16390), .CO(n16448), .S(n16393)
         );
  CMPR32X1 U4135 ( .A(n16580), .B(n16579), .C(n16578), .CO(n16711), .S(n16590)
         );
  CMPR32X1 U4136 ( .A(n7046), .B(n7045), .C(n7044), .CO(n7109), .S(n7082) );
  CMPR32X1 U4137 ( .A(n7031), .B(n7030), .C(n7029), .CO(n7081), .S(n7078) );
  CMPR32X1 U4138 ( .A(n6864), .B(n6865), .C(n6863), .CO(n6874), .S(n6853) );
  CMPR32X1 U4139 ( .A(n6973), .B(n6972), .C(n6971), .CO(n7080), .S(n6995) );
  CMPR32X1 U4140 ( .A(n9359), .B(n9545), .C(n9544), .CO(n9588), .S(n9539) );
  CMPR32X1 U4141 ( .A(n7101), .B(n7100), .C(n7099), .CO(n7136), .S(n7105) );
  ADDFX2 U4142 ( .A(n18534), .B(n18533), .CI(n18532), .CO(n18559), .S(n18555)
         );
  ADDFX2 U4143 ( .A(n16601), .B(n16600), .CI(n16599), .CO(n16669), .S(n16662)
         );
  OAI21XL U4144 ( .A0(n5455), .A1(n18659), .B0(n5928), .Y(n17758) );
  OAI2BB1X1 U4145 ( .A0N(n13612), .A1N(n13611), .B0(n5151), .Y(n13752) );
  CMPR32X1 U4146 ( .A(n13897), .B(n13896), .C(n13895), .CO(n13924), .S(n13870)
         );
  NAND2X1 U4147 ( .A(n5778), .B(n5776), .Y(n12452) );
  OAI2BB1X1 U4148 ( .A0N(n5876), .A1N(n18350), .B0(n5875), .Y(n18374) );
  OAI2BB1X1 U4149 ( .A0N(n3562), .A1N(n6974), .B0(n3560), .Y(n7079) );
  OAI21X1 U4150 ( .A0(n3595), .A1(n3594), .B0(n3593), .Y(n6416) );
  ADDFHX1 U4151 ( .A(n13454), .B(n13453), .CI(n13452), .CO(n13484), .S(n13457)
         );
  ADDFHX1 U4152 ( .A(n13686), .B(n13685), .CI(n13684), .CO(n13748), .S(n13753)
         );
  ADDFHX1 U4153 ( .A(n11742), .B(n11741), .CI(n11740), .CO(n11791), .S(n11827)
         );
  ADDFHX1 U4154 ( .A(n13559), .B(n13558), .CI(n13557), .CO(n13626), .S(n13585)
         );
  ADDFHX1 U4155 ( .A(n10418), .B(n10417), .CI(n10416), .CO(n10422), .S(n10435)
         );
  ADDFHX1 U4156 ( .A(n9638), .B(n9637), .CI(n9636), .CO(n10094), .S(n9662) );
  ADDFHX1 U4157 ( .A(n13304), .B(n13303), .CI(n13302), .CO(n13337), .S(n13305)
         );
  XNOR2X1 U4158 ( .A(n5304), .B(n9478), .Y(n5303) );
  ADDFHX1 U4159 ( .A(n12662), .B(n12661), .CI(n12660), .CO(n12667), .S(n12670)
         );
  ADDFHX1 U4160 ( .A(n13641), .B(n13640), .CI(n13639), .CO(n13811), .S(n13623)
         );
  CMPR32X1 U4161 ( .A(n12607), .B(n12606), .C(n12605), .CO(n12609), .S(n12666)
         );
  OAI21X2 U4162 ( .A0(n4070), .A1(n4349), .B0(n3281), .Y(n3280) );
  ADDFHX1 U4163 ( .A(n11841), .B(n11840), .CI(n11839), .CO(n11836), .S(n12432)
         );
  ADDFHX1 U4164 ( .A(n11705), .B(n11704), .CI(n11703), .CO(n11757), .S(n11713)
         );
  XOR3X2 U4165 ( .A(n16428), .B(n5802), .C(n16427), .Y(n16436) );
  ADDFHX2 U4166 ( .A(n17557), .B(n17556), .CI(n17555), .CO(n17627), .S(n17609)
         );
  ADDFHX2 U4167 ( .A(n6950), .B(n6949), .CI(n6948), .CO(n6982), .S(n6952) );
  CMPR32X1 U4168 ( .A(n18016), .B(n18015), .C(n18014), .CO(n18009), .S(n18098)
         );
  ADDFHX2 U4169 ( .A(n13480), .B(n13479), .CI(n13478), .CO(n13517), .S(n13502)
         );
  OAI21XL U4170 ( .A0(n13611), .A1(n13612), .B0(n13610), .Y(n5151) );
  ADDFHX2 U4171 ( .A(n7037), .B(n7036), .CI(n7035), .CO(n7085), .S(n7074) );
  CMPR32X1 U4172 ( .A(n12627), .B(n12626), .C(n12625), .CO(n12661), .S(n12665)
         );
  CMPR32X1 U4173 ( .A(n12538), .B(n12537), .C(n12536), .CO(n12552), .S(n12607)
         );
  ADDFX2 U4174 ( .A(n12048), .B(n12047), .CI(n12046), .CO(n12438), .S(n12455)
         );
  CMPR32X1 U4175 ( .A(n6740), .B(n6739), .C(n6738), .CO(n6764), .S(n6799) );
  CMPR32X1 U4176 ( .A(n6755), .B(n6754), .C(n6753), .CO(n6767), .S(n6795) );
  ADDFX2 U4177 ( .A(n18094), .B(n18093), .CI(n18092), .CO(n18076), .S(n18271)
         );
  CMPR32X1 U4178 ( .A(n15989), .B(n15988), .C(n15987), .CO(n16042), .S(n15994)
         );
  CMPR32X1 U4179 ( .A(n11679), .B(n11678), .C(n11677), .CO(n11682), .S(n11740)
         );
  CMPR32X1 U4180 ( .A(n13071), .B(n13070), .C(n13069), .CO(n13147), .S(n13146)
         );
  ADDFX2 U4181 ( .A(n6687), .B(n6686), .CI(n6685), .CO(n6702), .S(n6698) );
  CMPR32X1 U4182 ( .A(n18126), .B(n18125), .C(n18124), .CO(n18210), .S(n18209)
         );
  CMPR32X1 U4183 ( .A(n6339), .B(n6338), .C(n6337), .CO(n6800), .S(n6335) );
  CMPR32X1 U4184 ( .A(n12008), .B(n12007), .C(n12006), .CO(n12435), .S(n12451)
         );
  CMPR32X1 U4185 ( .A(n17661), .B(n17660), .C(n17659), .CO(n17667), .S(n17683)
         );
  ADDFX2 U4186 ( .A(n11669), .B(n11668), .CI(n11667), .CO(n11717), .S(n11680)
         );
  OAI21XL U4187 ( .A0(n4570), .A1(n9402), .B0(n3292), .Y(n9426) );
  OAI21XL U4188 ( .A0(n13649), .A1(n14249), .B0(n4933), .Y(n13689) );
  OAI21XL U4189 ( .A0(n3287), .A1(n9209), .B0(n3301), .Y(n9278) );
  OAI21XL U4190 ( .A0(n3940), .A1(n3466), .B0(n3464), .Y(n12094) );
  OAI21XL U4191 ( .A0(n3287), .A1(n10333), .B0(n3296), .Y(n10371) );
  CMPR32X1 U4192 ( .A(n12366), .B(n12365), .C(n12364), .CO(n12371), .S(n12373)
         );
  CMPR32X1 U4193 ( .A(n17618), .B(n17617), .C(n17616), .CO(n17769), .S(n17610)
         );
  CMPR32X1 U4194 ( .A(n6383), .B(n6382), .C(n6381), .CO(n6391), .S(n6421) );
  CMPR32X1 U4195 ( .A(n10342), .B(n10341), .C(n10340), .CO(n10359), .S(n10415)
         );
  CMPR32X1 U4196 ( .A(n6464), .B(n6463), .C(n6462), .CO(n6696), .S(n6676) );
  CMPR32X1 U4197 ( .A(n13969), .B(n13968), .C(n13967), .CO(n14036), .S(n13964)
         );
  OAI21XL U4198 ( .A0(n4570), .A1(n9230), .B0(n3289), .Y(n9246) );
  OAI21XL U4199 ( .A0(n3287), .A1(n9616), .B0(n3298), .Y(n9621) );
  OAI21XL U4200 ( .A0(n15979), .A1(n16688), .B0(n5759), .Y(n15978) );
  ADDFX2 U4201 ( .A(n9872), .B(n9871), .CI(n9870), .CO(n9944), .S(n9937) );
  CMPR32X1 U4202 ( .A(n11761), .B(n11760), .C(n11759), .CO(n11898), .S(n11753)
         );
  CMPR32X1 U4203 ( .A(n11632), .B(n11631), .C(n11630), .CO(n11755), .S(n11715)
         );
  ADDFX2 U4204 ( .A(n9620), .B(n9619), .CI(n9618), .CO(n10082), .S(n9648) );
  INVX1 U4205 ( .A(n5805), .Y(n5802) );
  OAI21XL U4206 ( .A0(n18541), .A1(n18538), .B0(n5895), .Y(n18550) );
  ADDFX2 U4207 ( .A(n16131), .B(n16130), .CI(n16129), .CO(n16160), .S(n16147)
         );
  ADDFX2 U4208 ( .A(n12564), .B(n12563), .CI(n12562), .CO(n12568), .S(n12547)
         );
  ADDFX2 U4209 ( .A(n9758), .B(n9757), .CI(n9756), .CO(n9770), .S(n9790) );
  ADDFX2 U4210 ( .A(n10365), .B(n10364), .CI(n10363), .CO(n10375), .S(n10358)
         );
  OAI2BB1X2 U4211 ( .A0N(n4066), .A1N(n17932), .B0(n4065), .Y(n18378) );
  OAI21XL U4212 ( .A0(n15592), .A1(n15598), .B0(n15593), .Y(n15629) );
  OAI21XL U4213 ( .A0(n15530), .A1(n15529), .B0(n15528), .Y(n15531) );
  OAI21XL U4214 ( .A0(n8781), .A1(n8780), .B0(n8779), .Y(n8782) );
  OAI2BB1X1 U4215 ( .A0N(n9796), .A1N(n5185), .B0(n5184), .Y(n9791) );
  OAI2BB1X1 U4216 ( .A0N(n3731), .A1N(n11665), .B0(n3730), .Y(n11716) );
  OAI21XL U4217 ( .A0(n3160), .A1(n8825), .B0(n8824), .Y(n8835) );
  OAI21XL U4218 ( .A0(n14967), .A1(n15575), .B0(n15574), .Y(n15585) );
  OAI21XL U4219 ( .A0(n8842), .A1(n8848), .B0(n8843), .Y(n8879) );
  ADDFHX1 U4220 ( .A(n17914), .B(n17913), .CI(n17912), .CO(n18379), .S(n17954)
         );
  ADDFHX1 U4221 ( .A(n17961), .B(n17960), .CI(n17959), .CO(n17953), .S(n17988)
         );
  ADDFHX1 U4222 ( .A(n12193), .B(n12192), .CI(n12191), .CO(n12216), .S(n12194)
         );
  OAI21XL U4223 ( .A0(n22030), .A1(n22036), .B0(n22031), .Y(n22067) );
  ADDFHX1 U4224 ( .A(n13236), .B(n13235), .CI(n13234), .CO(n13241), .S(n13243)
         );
  ADDFHX1 U4225 ( .A(n12057), .B(n12056), .CI(n12055), .CO(n12062), .S(n12089)
         );
  ADDFX2 U4226 ( .A(n17670), .B(n17669), .CI(n17668), .CO(n17665), .S(n18337)
         );
  NOR2X1 U4227 ( .A(n18740), .B(n4521), .Y(n19026) );
  ADDFHX1 U4228 ( .A(n17653), .B(n17652), .CI(n17651), .CO(n17608), .S(n17689)
         );
  ADDFHX1 U4229 ( .A(n6690), .B(n6689), .CI(n6688), .CO(n6697), .S(n6693) );
  ADDFX2 U4230 ( .A(n18260), .B(n18259), .CI(n18258), .CO(n18262), .S(n18211)
         );
  ADDFHX1 U4231 ( .A(n18288), .B(n18287), .CI(n18286), .CO(n18290), .S(n18265)
         );
  ADDFX2 U4232 ( .A(n9743), .B(n9742), .CI(n9741), .CO(n9738), .S(n9829) );
  CMPR32X1 U4233 ( .A(n17949), .B(n17948), .C(n17947), .CO(n17960), .S(n17989)
         );
  CMPR32X1 U4234 ( .A(n18276), .B(n18275), .C(n18274), .CO(n18092), .S(n18285)
         );
  CMPR32X1 U4235 ( .A(n13373), .B(n13374), .C(n13372), .CO(n13386), .S(n13370)
         );
  CMPR32X1 U4236 ( .A(n18251), .B(n18250), .C(n18249), .CO(n18256), .S(n18258)
         );
  CMPR32X1 U4237 ( .A(n12390), .B(n12389), .C(n12388), .CO(n12210), .S(n12399)
         );
  CMPR32X1 U4238 ( .A(n13232), .B(n13233), .C(n13231), .CO(n13299), .S(n13242)
         );
  CMPR32X1 U4239 ( .A(n13214), .B(n13213), .C(n13212), .CO(n13238), .S(n13234)
         );
  CMPR32X1 U4240 ( .A(n12000), .B(n11999), .C(n11998), .CO(n12448), .S(n12453)
         );
  CMPR32X1 U4241 ( .A(n12039), .B(n12038), .C(n12037), .CO(n12059), .S(n12055)
         );
  CMPR32X1 U4242 ( .A(n6786), .B(n6787), .C(n6785), .CO(n6792), .S(n6797) );
  OAI21XL U4243 ( .A0(n10328), .A1(n4570), .B0(n3290), .Y(n10351) );
  OAI2BB1X1 U4244 ( .A0N(n17546), .A1N(n17545), .B0(n5924), .Y(n17555) );
  CMPR32X1 U4245 ( .A(n16283), .B(n11953), .C(n11952), .CO(n11991), .S(n11947)
         );
  ADDFX2 U4246 ( .A(n13726), .B(n13725), .CI(n13724), .CO(n13783), .S(n13731)
         );
  CMPR32X1 U4247 ( .A(n12130), .B(n12129), .C(n12128), .CO(n12122), .S(n12160)
         );
  CMPR32X1 U4248 ( .A(n18062), .B(n18061), .C(n18060), .CO(n18074), .S(n18094)
         );
  ADDFX2 U4249 ( .A(n9661), .B(n9660), .CI(n9659), .CO(n9663), .S(n9690) );
  CMPR32X1 U4250 ( .A(n9752), .B(n9751), .C(n9750), .CO(n9747), .S(n9792) );
  CMPR32X1 U4251 ( .A(n13799), .B(n13798), .C(n13797), .CO(n13854), .S(n13785)
         );
  CMPR32X1 U4252 ( .A(n12259), .B(n12258), .C(n12257), .CO(n12252), .S(n12261)
         );
  CMPR32X1 U4253 ( .A(n12601), .B(n12600), .C(n12599), .CO(n12587), .S(n12625)
         );
  CMPR32X1 U4254 ( .A(n6818), .B(n6817), .C(n6816), .CO(n6880), .S(n6883) );
  ADDFX2 U4255 ( .A(n6536), .B(n4758), .CI(n6534), .CO(n6681), .S(n6532) );
  ADDFX2 U4256 ( .A(n17981), .B(n17980), .CI(n17979), .CO(n17991), .S(n18014)
         );
  INVX1 U4257 ( .A(n13665), .Y(n13602) );
  OAI21XL U4258 ( .A0(n12717), .A1(n11745), .B0(n5790), .Y(n5789) );
  OAI21XL U4259 ( .A0(n16049), .A1(n16704), .B0(n3698), .Y(n3697) );
  INVX1 U4260 ( .A(n11846), .Y(n4422) );
  ADDFX2 U4261 ( .A(n12363), .B(n12362), .CI(n12361), .CO(n12392), .S(n12372)
         );
  ADDFX2 U4262 ( .A(n9849), .B(n9848), .CI(n9847), .CO(n9990), .S(n9860) );
  ADDFX2 U4263 ( .A(n18091), .B(n18090), .CI(n18089), .CO(n18078), .S(n18280)
         );
  ADDFX2 U4264 ( .A(n6628), .B(n6627), .CI(n6626), .CO(n6630), .S(n6592) );
  XOR2X1 U4265 ( .A(n4356), .B(n10297), .Y(n10303) );
  OAI2BB1X1 U4266 ( .A0N(n4445), .A1N(n11729), .B0(n4444), .Y(n11739) );
  OAI21XL U4267 ( .A0(n3165), .A1(n19954), .B0(n19953), .Y(n19964) );
  OAI2BB1X1 U4268 ( .A0N(n6051), .A1N(n13732), .B0(n6050), .Y(n13786) );
  OAI22X2 U4269 ( .A0(n4570), .A1(n9361), .B0(n10403), .B1(n6139), .Y(n9478)
         );
  ADDFHX1 U4270 ( .A(n9705), .B(n9704), .CI(n9703), .CO(n9717), .S(n9739) );
  ADDFHX1 U4271 ( .A(n9727), .B(n9726), .CI(n9725), .CO(n9740), .S(n9760) );
  ADDFHX1 U4272 ( .A(n17891), .B(n17890), .CI(n17889), .CO(n18348), .S(n17913)
         );
  XNOR2X1 U4273 ( .A(n5372), .B(n3925), .Y(n3924) );
  ADDFHX1 U4274 ( .A(n13735), .B(n13734), .CI(n13733), .CO(n13787), .S(n13730)
         );
  ADDFX2 U4275 ( .A(n16016), .B(n16015), .CI(n16014), .CO(n16062), .S(n16099)
         );
  ADDFX2 U4276 ( .A(n17878), .B(n17877), .CI(n17876), .CO(n18364), .S(n18347)
         );
  CMPR32X1 U4277 ( .A(n9714), .B(n9713), .C(n9712), .CO(n9720), .S(n9741) );
  CMPR32X1 U4278 ( .A(n18116), .B(n18115), .C(n18114), .CO(n18249), .S(n18126)
         );
  CMPR32X1 U4279 ( .A(n12271), .B(n11658), .C(n17559), .CO(n17634), .S(n17561)
         );
  CMPR32X1 U4280 ( .A(n18031), .B(n18030), .C(n18029), .CO(n18040), .S(n18057)
         );
  OAI21XL U4281 ( .A0(n12995), .A1(n3110), .B0(n12535), .Y(n11676) );
  ADDFX2 U4282 ( .A(n11857), .B(n11856), .CI(n11855), .CO(n12445), .S(n12433)
         );
  CLKBUFX8 U4283 ( .A(n17087), .Y(n17074) );
  ADDFX2 U4284 ( .A(n12209), .B(n12208), .CI(n12207), .CO(n12197), .S(n12394)
         );
  ADDFX2 U4285 ( .A(n3049), .B(n3197), .CI(n11986), .CO(n12624), .S(n11981) );
  BUFX4 U4286 ( .A(n16330), .Y(n3102) );
  ADDFX2 U4287 ( .A(n18233), .B(n18232), .CI(n18231), .CO(n18279), .S(n18253)
         );
  ADDFX2 U4288 ( .A(n17917), .B(n17916), .CI(n17915), .CO(n18370), .S(n17933)
         );
  INVX1 U4289 ( .A(M0_b_1_), .Y(n7056) );
  OAI21XL U4290 ( .A0(n19910), .A1(n19909), .B0(n19908), .Y(n19911) );
  XOR2X1 U4291 ( .A(n4492), .B(n4490), .Y(n3870) );
  OAI21XL U4292 ( .A0(n3160), .A1(n8807), .B0(n8806), .Y(n8821) );
  OAI21XL U4293 ( .A0(n14967), .A1(n15556), .B0(n15555), .Y(n15571) );
  OAI21XL U4294 ( .A0(n3160), .A1(n8792), .B0(n8791), .Y(n8813) );
  OAI21XL U4295 ( .A0(n21854), .A1(n21996), .B0(n21995), .Y(n22010) );
  OAI21XL U4296 ( .A0(n14967), .A1(n15551), .B0(n15550), .Y(n15567) );
  OAI21XL U4297 ( .A0(n21854), .A1(n21991), .B0(n21990), .Y(n22006) );
  OAI21XL U4298 ( .A0(n14967), .A1(n15541), .B0(n15540), .Y(n15563) );
  OAI21XL U4299 ( .A0(n3160), .A1(n8797), .B0(n8796), .Y(n8815) );
  OAI21XL U4300 ( .A0(n14967), .A1(n15546), .B0(n15545), .Y(n15565) );
  OAI21XL U4301 ( .A0(n3160), .A1(n8787), .B0(n8786), .Y(n8811) );
  OAI21XL U4302 ( .A0(n21854), .A1(n21976), .B0(n21975), .Y(n22000) );
  NAND2X4 U4303 ( .A(n17061), .B(n3395), .Y(n17060) );
  XNOR2X1 U4304 ( .A(n10170), .B(n5541), .Y(n10167) );
  OAI21XL U4305 ( .A0(n19971), .A1(n19977), .B0(n19972), .Y(n20008) );
  NOR2X1 U4306 ( .A(n4425), .B(n4424), .Y(n4423) );
  OAI21X1 U4307 ( .A0(n3287), .A1(n9579), .B0(n3295), .Y(n10165) );
  OAI21XL U4308 ( .A0(n21838), .A1(n21947), .B0(n21837), .Y(n21972) );
  ADDFHX1 U4309 ( .A(n17998), .B(n17997), .CI(n17996), .CO(n18010), .S(n18033)
         );
  ADDFHX1 U4310 ( .A(n9733), .B(n9732), .CI(n9731), .CO(n9725), .S(n9769) );
  ADDFX2 U4311 ( .A(n9698), .B(n9697), .CI(n9696), .CO(n9705), .S(n9726) );
  CLKBUFX3 U4312 ( .A(n16570), .Y(n16701) );
  BUFX3 U4313 ( .A(n17073), .Y(n5677) );
  ADDFHX2 U4314 ( .A(n17978), .B(n17977), .CI(n17976), .CO(n17971), .S(n18015)
         );
  CLKINVX3 U4315 ( .A(n6347), .Y(n7634) );
  BUFX3 U4316 ( .A(n17147), .Y(n3194) );
  OAI21XL U4317 ( .A0(n4570), .A1(n9549), .B0(n3291), .Y(n9585) );
  OAI21XL U4318 ( .A0(n11794), .A1(n12284), .B0(n3918), .Y(n3917) );
  INVX4 U4319 ( .A(n16572), .Y(n16289) );
  BUFX3 U4320 ( .A(n16686), .Y(n16638) );
  INVX4 U4321 ( .A(n6744), .Y(n7712) );
  BUFX3 U4322 ( .A(n15947), .Y(n16699) );
  OAI2BB1X1 U4323 ( .A0N(n13899), .A1N(n2997), .B0(n13898), .Y(n13928) );
  BUFX4 U4324 ( .A(n16867), .Y(n16941) );
  BUFX3 U4325 ( .A(n15949), .Y(n16939) );
  OAI21XL U4326 ( .A0(n3165), .A1(n19931), .B0(n19930), .Y(n19946) );
  OAI21XL U4327 ( .A0(n3165), .A1(n19926), .B0(n19925), .Y(n19944) );
  INVX1 U4328 ( .A(n3686), .Y(n3018) );
  BUFX4 U4329 ( .A(n10532), .Y(n10517) );
  NAND2X1 U4330 ( .A(n16319), .B(n5096), .Y(n17087) );
  OAI21X2 U4331 ( .A0(n3287), .A1(n9701), .B0(n3293), .Y(n9732) );
  AOI2BB1X1 U4332 ( .A0N(n18659), .A1N(n17672), .B0(n4491), .Y(n4490) );
  INVX1 U4333 ( .A(n5835), .Y(n3044) );
  BUFX3 U4334 ( .A(n10329), .Y(n3174) );
  XOR2X1 U4335 ( .A(n5543), .B(n5542), .Y(n5541) );
  ADDFHX1 U4336 ( .A(n17532), .B(n17531), .CI(n17530), .CO(n17576), .S(n17545)
         );
  CLKINVX3 U4337 ( .A(n3213), .Y(n7286) );
  INVX4 U4338 ( .A(n17038), .Y(n17039) );
  BUFX3 U4339 ( .A(n12746), .Y(n12525) );
  BUFX3 U4340 ( .A(n10369), .Y(n9780) );
  INVX4 U4341 ( .A(n10540), .Y(n25885) );
  CLKBUFX3 U4342 ( .A(M2_b_19_), .Y(n10538) );
  OAI21XL U4343 ( .A0(n3287), .A1(n9666), .B0(n3300), .Y(n9677) );
  INVX4 U4344 ( .A(n5079), .Y(n10494) );
  OAI21XL U4345 ( .A0(n17604), .A1(n18226), .B0(n6034), .Y(n17607) );
  BUFX4 U4346 ( .A(n9590), .Y(n9979) );
  OAI21XL U4347 ( .A0(n3160), .A1(n8771), .B0(n8770), .Y(n8776) );
  OAI21XL U4348 ( .A0(n14967), .A1(n15520), .B0(n15519), .Y(n15525) );
  BUFX3 U4349 ( .A(n9215), .Y(n10533) );
  OAI2BB1X1 U4350 ( .A0N(n12107), .A1N(n5981), .B0(n5979), .Y(n3939) );
  INVX1 U4351 ( .A(n6300), .Y(n6347) );
  INVX1 U4352 ( .A(n10171), .Y(n5542) );
  AOI21X1 U4353 ( .A0(n4915), .A1(n4916), .B0(n4889), .Y(n4914) );
  ADDFX2 U4354 ( .A(n4750), .B(n17584), .CI(n17583), .CO(n17594), .S(n17666)
         );
  BUFX3 U4355 ( .A(M2_b_18_), .Y(n10539) );
  BUFX3 U4356 ( .A(M2_b_7_), .Y(n9839) );
  BUFX4 U4357 ( .A(n15996), .Y(n3105) );
  CLKINVX3 U4358 ( .A(n6366), .Y(n6990) );
  CLKBUFX8 U4359 ( .A(n16893), .Y(n16977) );
  CLKBUFX3 U4360 ( .A(M2_b_6_), .Y(n9836) );
  INVX4 U4361 ( .A(n10338), .Y(n10339) );
  INVX4 U4362 ( .A(n13173), .Y(n3173) );
  OAI21XL U4363 ( .A0(n12597), .A1(n12126), .B0(n6102), .Y(n12142) );
  OAI21XL U4364 ( .A0(n9652), .A1(n10496), .B0(n5149), .Y(n5148) );
  CLKINVX3 U4365 ( .A(n5298), .Y(n10540) );
  CLKBUFX8 U4366 ( .A(n4570), .Y(n3287) );
  CLKINVX3 U4367 ( .A(n5087), .Y(n5086) );
  CLKBUFX8 U4368 ( .A(M0_b_17_), .Y(n7646) );
  BUFX3 U4369 ( .A(M2_b_12_), .Y(n10387) );
  BUFX4 U4370 ( .A(n12521), .Y(n12995) );
  INVX1 U4371 ( .A(n4797), .Y(n3200) );
  INVX1 U4372 ( .A(n3196), .Y(n5997) );
  NAND2X4 U4373 ( .A(n11625), .B(n12070), .Y(n12152) );
  INVX1 U4374 ( .A(n5399), .Y(n5398) );
  NAND2X1 U4375 ( .A(n4532), .B(n4529), .Y(M5_a_6_) );
  INVX1 U4376 ( .A(n6291), .Y(n7534) );
  BUFX4 U4377 ( .A(n9781), .Y(n3180) );
  INVX4 U4378 ( .A(n7564), .Y(n25869) );
  INVX1 U4379 ( .A(n14291), .Y(n13510) );
  INVX1 U4380 ( .A(n3288), .Y(n3297) );
  BUFX3 U4381 ( .A(M2_b_13_), .Y(n10386) );
  OAI21XL U4382 ( .A0(n15400), .A1(n15507), .B0(n15399), .Y(n15532) );
  INVX1 U4383 ( .A(M5_mult_x_15_n1), .Y(n3205) );
  XNOR2X1 U4384 ( .A(M2_a_12_), .B(n10338), .Y(n9203) );
  NAND3X1 U4385 ( .A(n6019), .B(n6020), .C(n6018), .Y(M5_a_22_) );
  XNOR2X1 U4386 ( .A(n6291), .B(n5399), .Y(n6326) );
  BUFX3 U4387 ( .A(n25243), .Y(n3115) );
  XOR2X2 U4388 ( .A(M0_a_22_), .B(n6746), .Y(n7826) );
  BUFX8 U4389 ( .A(n4569), .Y(n4570) );
  CLKBUFX3 U4390 ( .A(M0_b_7_), .Y(n25881) );
  BUFX3 U4391 ( .A(M0_b_4_), .Y(n7165) );
  INVX4 U4392 ( .A(n3210), .Y(n18453) );
  CLKBUFX3 U4393 ( .A(M2_b_2_), .Y(n9892) );
  INVX4 U4394 ( .A(n6829), .Y(n25867) );
  CLKINVX3 U4395 ( .A(M3_mult_x_15_n1682), .Y(n16965) );
  OAI21XL U4396 ( .A0(n12618), .A1(n11957), .B0(n5940), .Y(n5939) );
  BUFX3 U4397 ( .A(n15970), .Y(M5_mult_x_15_n1) );
  CLKBUFX8 U4398 ( .A(n12578), .Y(n12717) );
  CLKINVX3 U4399 ( .A(M2_a_19_), .Y(n5079) );
  INVX4 U4400 ( .A(n6989), .Y(n25866) );
  INVX1 U4401 ( .A(n18503), .Y(n3189) );
  INVX1 U4402 ( .A(M3_mult_x_15_b_19_), .Y(n5718) );
  OAI2BB1X1 U4403 ( .A0N(n6035), .A1N(n3192), .B0(n3392), .Y(n17589) );
  INVXL U4404 ( .A(n5646), .Y(n5645) );
  INVX1 U4405 ( .A(n4783), .Y(n4784) );
  BUFX3 U4406 ( .A(n12070), .Y(n3185) );
  OAI21XL U4407 ( .A0(n25243), .A1(n26234), .B0(n11523), .Y(M1_a_11_) );
  OAI21XL U4408 ( .A0(n25243), .A1(n25901), .B0(n11524), .Y(M1_a_12_) );
  BUFX4 U4409 ( .A(M2_b_4_), .Y(n9874) );
  NAND2X1 U4410 ( .A(n5448), .B(n5447), .Y(n5811) );
  NAND2BX1 U4411 ( .AN(n4534), .B(n4533), .Y(M5_a_10_) );
  INVX1 U4412 ( .A(n13899), .Y(n13057) );
  XOR2X1 U4413 ( .A(M0_a_6_), .B(n7092), .Y(n5583) );
  INVX2 U4414 ( .A(n6746), .Y(n7711) );
  INVX1 U4415 ( .A(n4794), .Y(n4795) );
  BUFX3 U4416 ( .A(n11749), .Y(n12760) );
  NAND3BX1 U4417 ( .AN(n5080), .B(n9082), .C(n9081), .Y(n5255) );
  NOR2X2 U4418 ( .A(n3476), .B(n3475), .Y(n5399) );
  INVX1 U4419 ( .A(n13898), .Y(n13842) );
  NAND2X1 U4420 ( .A(n4558), .B(n3478), .Y(n6291) );
  AOI2BB2X1 U4421 ( .B0(n3383), .B1(n3382), .A0N(n3183), .A1N(n3941), .Y(n3846) );
  XOR2XL U4422 ( .A(n14228), .B(n5391), .Y(n13357) );
  NAND3BX1 U4423 ( .AN(n5204), .B(n9070), .C(n9069), .Y(M2_a_18_) );
  NAND3BX1 U4424 ( .AN(n24024), .B(n5608), .C(n5607), .Y(M0_a_22_) );
  XOR2XL U4425 ( .A(n6829), .B(n5628), .Y(n5627) );
  XOR2X1 U4426 ( .A(n6989), .B(n3591), .Y(n3590) );
  INVX1 U4427 ( .A(M1_b_19_), .Y(n14267) );
  XNOR2XL U4428 ( .A(n4945), .B(n4919), .Y(n11627) );
  BUFX4 U4429 ( .A(M2_b_10_), .Y(n10342) );
  NAND3BX1 U4430 ( .AN(n5492), .B(n9090), .C(n5491), .Y(M2_b_12_) );
  AOI2BB1X2 U4431 ( .A0N(n25767), .A1N(n26024), .B0(n5088), .Y(n5087) );
  NOR2X1 U4432 ( .A(n25767), .B(n26246), .Y(n3396) );
  BUFX3 U4433 ( .A(n11485), .Y(n12233) );
  BUFX8 U4434 ( .A(M3_mult_x_15_b_3_), .Y(n12279) );
  BUFX8 U4435 ( .A(M5_b_18_), .Y(n3196) );
  BUFX3 U4436 ( .A(n17605), .Y(n17832) );
  INVX4 U4437 ( .A(n9843), .Y(n9841) );
  BUFX8 U4438 ( .A(M3_mult_x_15_b_19_), .Y(n3048) );
  INVX4 U4439 ( .A(n18142), .Y(n18150) );
  CLKBUFX8 U4440 ( .A(M3_mult_x_15_n1682), .Y(n5430) );
  CLKINVX3 U4441 ( .A(M3_mult_x_15_b_20_), .Y(n4206) );
  CLKBUFX8 U4442 ( .A(M3_mult_x_15_b_21_), .Y(n12803) );
  INVX1 U4443 ( .A(M5_a_20_), .Y(n4794) );
  OAI211X4 U4444 ( .A0(n23998), .A1(n25243), .B0(n9102), .C0(n11508), .Y(
        M2_b_4_) );
  BUFX12 U4445 ( .A(M3_mult_x_15_b_6_), .Y(n3049) );
  CLKINVX3 U4446 ( .A(M0_a_7_), .Y(n6829) );
  CLKINVX4 U4447 ( .A(n5029), .Y(n18721) );
  CLKINVX3 U4448 ( .A(M3_a_22_), .Y(n3112) );
  CLKINVX3 U4449 ( .A(n17073), .Y(n3212) );
  OAI21XL U4450 ( .A0(n25243), .A1(n23993), .B0(n13040), .Y(n4322) );
  AND2X2 U4451 ( .A(n9083), .B(n4464), .Y(M2_U4_U1_or2_inv_0__26_) );
  NAND2X4 U4452 ( .A(n17494), .B(n18653), .Y(n18652) );
  OAI21XL U4453 ( .A0(n25243), .A1(n25907), .B0(n11518), .Y(M1_a_3_) );
  OAI21XL U4454 ( .A0(n25243), .A1(n25900), .B0(n11513), .Y(M1_a_2_) );
  BUFX3 U4455 ( .A(n18666), .Y(n18659) );
  XOR2X1 U4456 ( .A(n11480), .B(n3638), .Y(n12070) );
  NAND3BX2 U4457 ( .AN(n25158), .B(n5606), .C(n5605), .Y(n6746) );
  OAI21X2 U4458 ( .A0(n26030), .A1(n25767), .B0(n5647), .Y(n5646) );
  NAND2X1 U4459 ( .A(n11544), .B(n11543), .Y(M1_b_20_) );
  AOI2BB1X2 U4460 ( .A0N(n25796), .A1N(n26245), .B0(n5651), .Y(n16909) );
  XOR2XL U4461 ( .A(n4002), .B(n3638), .Y(n11625) );
  XNOR2X1 U4462 ( .A(n5045), .B(M3_U3_U1_or2_inv_0__18_), .Y(n4054) );
  XNOR2X1 U4463 ( .A(M0_a_8_), .B(M0_a_7_), .Y(n6294) );
  OAI21X2 U4464 ( .A0(n15941), .A1(n26270), .B0(n3678), .Y(n15970) );
  OAI21X2 U4465 ( .A0(n15941), .A1(n26295), .B0(n3676), .Y(M5_a_2_) );
  NOR2BX2 U4466 ( .AN(n9096), .B(n4250), .Y(n6076) );
  NAND2XL U4467 ( .A(n7389), .B(y10[22]), .Y(n5608) );
  NAND2BX1 U4468 ( .AN(n25152), .B(n3477), .Y(n3476) );
  NAND2X1 U4469 ( .A(n9164), .B(target_temp[21]), .Y(n13507) );
  OAI211X1 U4470 ( .A0(n23994), .A1(n25243), .B0(n9077), .C0(n11505), .Y(
        M2_b_8_) );
  NAND3X1 U4471 ( .A(n4662), .B(n5133), .C(n5132), .Y(M0_b_18_) );
  OAI211X1 U4472 ( .A0(n23989), .A1(n25243), .B0(n9100), .C0(n13356), .Y(
        M2_b_17_) );
  AOI21X1 U4473 ( .A0(n25206), .A1(data[103]), .B0(n3804), .Y(n3803) );
  OAI222X1 U4474 ( .A0(n26275), .A1(n4860), .B0(n25928), .B1(n25767), .C0(
        n26035), .C1(n15940), .Y(M5_a_18_) );
  XNOR2X2 U4475 ( .A(M1_b_18_), .B(n3019), .Y(n13428) );
  CLKBUFX3 U4476 ( .A(n12293), .Y(n12340) );
  OAI211X4 U4477 ( .A0(n25904), .A1(n9087), .B0(n9092), .C0(n9091), .Y(M2_a_8_) );
  BUFX4 U4478 ( .A(M2_b_0_), .Y(n9960) );
  CLKBUFX8 U4479 ( .A(M3_mult_x_15_b_14_), .Y(n18611) );
  CLKBUFX8 U4480 ( .A(n11498), .Y(M3_mult_x_15_b_3_) );
  CLKINVX3 U4481 ( .A(n14228), .Y(n3019) );
  AND2X2 U4482 ( .A(n18658), .B(n5470), .Y(n5029) );
  CLKBUFX8 U4483 ( .A(n12025), .Y(n12357) );
  INVXL U4484 ( .A(M4_a_12_), .Y(n5462) );
  NAND2X4 U4485 ( .A(n10496), .B(n5238), .Y(n9504) );
  INVX1 U4486 ( .A(n5045), .Y(n5044) );
  XOR2X1 U4487 ( .A(n4189), .B(n5374), .Y(n4396) );
  AND2X2 U4488 ( .A(n5262), .B(n11531), .Y(n3331) );
  NAND2X1 U4489 ( .A(n17495), .B(n17605), .Y(n18666) );
  INVX1 U4490 ( .A(n4434), .Y(n3740) );
  OAI21X2 U4491 ( .A0(n7382), .A1(n25995), .B0(n6226), .Y(M0_a_10_) );
  INVXL U4492 ( .A(n25158), .Y(n4340) );
  NAND3X1 U4493 ( .A(n9085), .B(n9084), .C(n5180), .Y(M2_a_10_) );
  NAND2X2 U4494 ( .A(n11527), .B(n11528), .Y(M1_b_15_) );
  OAI21XL U4495 ( .A0(n19781), .A1(n19887), .B0(n19780), .Y(n19912) );
  XNOR2XL U4496 ( .A(M3_mult_x_15_a_15_), .B(n4979), .Y(n5942) );
  NAND2X1 U4497 ( .A(n11534), .B(n11533), .Y(n5391) );
  NOR2X1 U4498 ( .A(n5649), .B(n5648), .Y(n5647) );
  NAND2BXL U4499 ( .AN(n9087), .B(n4720), .Y(n4341) );
  NAND2XL U4500 ( .A(n9164), .B(target_temp[19]), .Y(n11541) );
  NOR2XL U4501 ( .A(n25153), .B(n3574), .Y(n6259) );
  AOI21X2 U4502 ( .A0(sigma10[9]), .A1(n25206), .B0(n3333), .Y(n6162) );
  NOR2XL U4503 ( .A(n15940), .B(n25919), .Y(n3804) );
  NAND2XL U4504 ( .A(n4566), .B(learning_rate[7]), .Y(n5295) );
  OAI21X1 U4505 ( .A0(n6266), .A1(n26215), .B0(n5567), .Y(n5566) );
  XNOR2X2 U4506 ( .A(M4_a_9_), .B(n4189), .Y(n18501) );
  AOI21X1 U4507 ( .A0(n6733), .A1(y10[5]), .B0(n25143), .Y(n6243) );
  OAI21X1 U4508 ( .A0(n26264), .A1(n25796), .B0(n4048), .Y(M3_a_22_) );
  AOI21XL U4509 ( .A0(n11479), .A1(data[117]), .B0(n6016), .Y(n6015) );
  INVX4 U4510 ( .A(n3191), .Y(n25884) );
  INVX4 U4511 ( .A(n12225), .Y(n3204) );
  BUFX8 U4512 ( .A(M3_mult_x_15_b_15_), .Y(n3198) );
  BUFX16 U4513 ( .A(M3_mult_x_15_b_12_), .Y(n12561) );
  CLKBUFX8 U4514 ( .A(n2974), .Y(n3108) );
  BUFX3 U4515 ( .A(n11480), .Y(n12282) );
  NAND2X1 U4516 ( .A(n5375), .B(n5881), .Y(M4_a_4_) );
  NOR2BX1 U4517 ( .AN(n4897), .B(n3741), .Y(n4434) );
  NAND2X1 U4518 ( .A(n4540), .B(n4537), .Y(M3_a_20_) );
  NAND2X1 U4519 ( .A(n11521), .B(n11520), .Y(M1_b_10_) );
  NAND3X1 U4520 ( .A(n9202), .B(n5567), .C(n5181), .Y(n21055) );
  INVX1 U4521 ( .A(M4_a_19_), .Y(n18637) );
  OAI2BB1X1 U4522 ( .A0N(n5032), .A1N(data[78]), .B0(n17473), .Y(n4888) );
  NAND2X2 U4523 ( .A(n3229), .B(data_point[19]), .Y(n9071) );
  NOR2X1 U4524 ( .A(n4582), .B(n5008), .Y(n25158) );
  XNOR2X1 U4525 ( .A(M3_mult_x_15_a_15_), .B(M3_a_16_), .Y(n11628) );
  CLKBUFX8 U4526 ( .A(n11495), .Y(n3021) );
  NOR2BX1 U4527 ( .AN(n17478), .B(n4226), .Y(n5470) );
  CLKINVX3 U4528 ( .A(M4_a_13_), .Y(n3210) );
  NOR2X1 U4529 ( .A(n15940), .B(n25924), .Y(n6016) );
  NAND2XL U4530 ( .A(n25206), .B(n3003), .Y(n4535) );
  XNOR2X2 U4531 ( .A(n4979), .B(M3_U3_U1_or2_inv_0__18_), .Y(n12616) );
  XNOR2X2 U4532 ( .A(M4_a_17_), .B(M4_a_18_), .Y(n18653) );
  XNOR2X2 U4533 ( .A(M4_a_5_), .B(M4_a_6_), .Y(n17902) );
  OAI2BB1X1 U4534 ( .A0N(n3758), .A1N(data[36]), .B0(n4899), .Y(n3639) );
  NOR2XL U4535 ( .A(in_valid_d), .B(n3573), .Y(n3574) );
  BUFX2 U4536 ( .A(n11489), .Y(M3_mult_x_15_b_7_) );
  NOR2BX2 U4537 ( .AN(n5049), .B(n3231), .Y(n3376) );
  CLKINVX3 U4538 ( .A(M3_mult_x_15_a_15_), .Y(n3191) );
  AND2X2 U4539 ( .A(n5491), .B(n5342), .Y(n4272) );
  INVX2 U4540 ( .A(n18222), .Y(n2977) );
  XOR2X1 U4541 ( .A(M4_a_17_), .B(n3756), .Y(n4511) );
  BUFX4 U4542 ( .A(M3_mult_x_15_b_2_), .Y(n12271) );
  OAI21X2 U4543 ( .A0(n15941), .A1(n6213), .B0(n4038), .Y(M3_mult_x_15_b_11_)
         );
  NAND2X1 U4544 ( .A(n5504), .B(n6086), .Y(n5511) );
  NOR2XL U4545 ( .A(n15942), .B(n26517), .Y(n3782) );
  NAND2XL U4546 ( .A(n25206), .B(data[52]), .Y(n4540) );
  NOR2X1 U4547 ( .A(n5435), .B(n5433), .Y(n5432) );
  NAND2X1 U4548 ( .A(n5434), .B(n4722), .Y(n5431) );
  OAI22X2 U4549 ( .A0(n25796), .A1(n26244), .B0(n26007), .B1(n15940), .Y(n3783) );
  OAI22X2 U4550 ( .A0(n25813), .A1(n25927), .B0(n26273), .B1(n17167), .Y(n3625) );
  OAI21X1 U4551 ( .A0(n3103), .A1(n26235), .B0(n9047), .Y(n3307) );
  CLKINVX3 U4552 ( .A(n21628), .Y(n3042) );
  NAND2X1 U4553 ( .A(n4520), .B(n6089), .Y(n4196) );
  OAI21X2 U4554 ( .A0(n15941), .A1(n25908), .B0(n3879), .Y(M3_mult_x_15_a_15_)
         );
  INVX2 U4555 ( .A(M3_mult_x_15_b_5_), .Y(n2973) );
  NOR2X1 U4556 ( .A(n6258), .B(n4581), .Y(n25152) );
  NAND2X1 U4557 ( .A(n25206), .B(sigma10[11]), .Y(n4038) );
  NOR2X2 U4558 ( .A(n25813), .B(n2989), .Y(n4224) );
  NOR2X1 U4559 ( .A(n6246), .B(n4583), .Y(n25145) );
  NOR2X1 U4560 ( .A(n25767), .B(n26250), .Y(n3232) );
  OAI21X1 U4561 ( .A0(n4860), .A1(n26235), .B0(n4601), .Y(n4319) );
  NAND2X1 U4562 ( .A(n9164), .B(y12[9]), .Y(n3286) );
  NAND2BX1 U4563 ( .AN(n3438), .B(n2995), .Y(n18222) );
  NOR2X1 U4564 ( .A(n25767), .B(n26259), .Y(n3893) );
  NOR2X1 U4565 ( .A(n6285), .B(n4581), .Y(n25151) );
  AOI2BB1X2 U4566 ( .A0N(n25796), .A1N(n26240), .B0(n5971), .Y(n5983) );
  AOI21X1 U4567 ( .A0(target_temp[2]), .A1(n21166), .B0(n6155), .Y(n6023) );
  NOR2X1 U4568 ( .A(n5943), .B(n3880), .Y(n3879) );
  NAND2BX1 U4569 ( .AN(n4418), .B(n4417), .Y(M3_mult_x_15_b_5_) );
  INVXL U4570 ( .A(data_point[11]), .Y(n6224) );
  OAI21XL U4571 ( .A0(n15942), .A1(n4725), .B0(n4669), .Y(n4085) );
  OAI21XL U4572 ( .A0(n15942), .A1(n6179), .B0(n6010), .Y(n4418) );
  INVX1 U4573 ( .A(n17474), .Y(n3435) );
  NAND2X1 U4574 ( .A(n22227), .B(n21442), .Y(n21737) );
  NAND2X1 U4575 ( .A(n25206), .B(n4729), .Y(n4417) );
  NOR2X1 U4576 ( .A(n4581), .B(n3538), .Y(n25153) );
  CLKINVX4 U4577 ( .A(n6169), .Y(n3155) );
  OAI21XL U4578 ( .A0(n25992), .A1(n21329), .B0(n21443), .Y(n23115) );
  OR2X2 U4579 ( .A(n8598), .B(n9027), .Y(n6169) );
  INVXL U4580 ( .A(data_point[15]), .Y(n3538) );
  BUFX8 U4581 ( .A(n11483), .Y(n4860) );
  CLKINVX3 U4582 ( .A(n8823), .Y(n9027) );
  CLKINVX4 U4583 ( .A(n15363), .Y(n15573) );
  NOR2X1 U4584 ( .A(n8179), .B(n23761), .Y(n20377) );
  OR2X2 U4585 ( .A(n15345), .B(n23955), .Y(n14967) );
  INVX4 U4586 ( .A(n8601), .Y(n3154) );
  CLKINVX3 U4587 ( .A(n8537), .Y(n8601) );
  OAI21XL U4588 ( .A0(n21628), .A1(n21579), .B0(n21555), .Y(n21697) );
  NAND2XL U4589 ( .A(n15792), .B(n14962), .Y(n15345) );
  NOR2X1 U4590 ( .A(n8178), .B(n8177), .Y(n20378) );
  CLKINVX3 U4591 ( .A(n6192), .Y(n3164) );
  OAI21XL U4592 ( .A0(n19237), .A1(n26227), .B0(n14963), .Y(n23170) );
  OR2X2 U4593 ( .A(n19683), .B(n3215), .Y(n6192) );
  OAI21XL U4594 ( .A0(n3040), .A1(n7890), .B0(n8194), .Y(n23178) );
  NOR2X1 U4595 ( .A(n20137), .B(n19345), .Y(n19683) );
  OAI21XL U4596 ( .A0(n3040), .A1(n8191), .B0(n8190), .Y(n23179) );
  OAI21XL U4597 ( .A0(n21519), .A1(n21408), .B0(n21407), .Y(n23121) );
  NOR2X1 U4598 ( .A(n19309), .B(n24310), .Y(n20137) );
  OAI21XL U4599 ( .A0(n3063), .A1(n26195), .B0(n19347), .Y(n23202) );
  OAI21XL U4600 ( .A0(n8228), .A1(n8231), .B0(n8229), .Y(n8272) );
  OAI21XL U4601 ( .A0(n3040), .A1(n8187), .B0(n8186), .Y(n23180) );
  OAI21XL U4602 ( .A0(n3040), .A1(n8183), .B0(n8182), .Y(n23181) );
  INVX1 U4603 ( .A(n24309), .Y(n24310) );
  BUFX3 U4604 ( .A(n15128), .Y(n15055) );
  CLKINVX3 U4605 ( .A(n4457), .Y(n6194) );
  OAI21XL U4606 ( .A0(n3020), .A1(n21433), .B0(n21432), .Y(n23123) );
  OAI21XL U4607 ( .A0(n3020), .A1(n21437), .B0(n21436), .Y(n23122) );
  CLKINVX3 U4608 ( .A(n19542), .Y(n3036) );
  INVX4 U4609 ( .A(n2996), .Y(n19807) );
  OAI21XL U4610 ( .A0(n3040), .A1(n8210), .B0(n8209), .Y(n23182) );
  CLKINVX3 U4611 ( .A(n8259), .Y(n8592) );
  OAI21XL U4612 ( .A0(n3040), .A1(n8206), .B0(n8205), .Y(n23183) );
  INVX1 U4613 ( .A(n4790), .Y(n4791) );
  INVX1 U4614 ( .A(n4792), .Y(n4793) );
  INVX4 U4615 ( .A(n15289), .Y(n3038) );
  OAI21XL U4616 ( .A0(n15558), .A1(n14929), .B0(n14928), .Y(n23160) );
  OAI21XL U4617 ( .A0(n3040), .A1(n8202), .B0(n8201), .Y(n23184) );
  OAI21XL U4618 ( .A0(n19564), .A1(n19317), .B0(n19316), .Y(n23205) );
  INVX1 U4619 ( .A(n4786), .Y(n4787) );
  OAI21XL U4620 ( .A0(n15558), .A1(n14957), .B0(n14956), .Y(n23161) );
  CLKINVX3 U4621 ( .A(n19510), .Y(n3094) );
  OAI21XL U4622 ( .A0(n3041), .A1(n19340), .B0(n19339), .Y(n23207) );
  OAI21XL U4623 ( .A0(n15558), .A1(n14953), .B0(n14952), .Y(n23162) );
  OAI21XL U4624 ( .A0(n3041), .A1(n19336), .B0(n19335), .Y(n23208) );
  CLKINVX3 U4625 ( .A(n19297), .Y(n19566) );
  OAI21XL U4626 ( .A0(n8023), .A1(n8022), .B0(n8021), .Y(n8024) );
  OAI21XL U4627 ( .A0(n8134), .A1(n8133), .B0(n8132), .Y(n8157) );
  OAI21XL U4628 ( .A0(n6173), .A1(n21311), .B0(n21328), .Y(n21417) );
  OAI21XL U4629 ( .A0(n6167), .A1(n21333), .B0(n21306), .Y(n21421) );
  OAI21XL U4630 ( .A0(n26159), .A1(n21329), .B0(n21327), .Y(n21418) );
  OAI21XL U4631 ( .A0(n19237), .A1(n7884), .B0(n7883), .Y(n8192) );
  OAI21XL U4632 ( .A0(n14901), .A1(n14900), .B0(n14899), .Y(n14902) );
  INVX1 U4633 ( .A(n8193), .Y(n8148) );
  OAI21XL U4634 ( .A0(n14833), .A1(n26546), .B0(n8096), .Y(n8207) );
  OAI21XL U4635 ( .A0(n19237), .A1(n8066), .B0(n8065), .Y(n8195) );
  OAI21XL U4636 ( .A0(n14813), .A1(n14812), .B0(n14811), .Y(n14814) );
  OAI21XL U4637 ( .A0(n14833), .A1(n26594), .B0(n8109), .Y(n8188) );
  OAI21XL U4638 ( .A0(n19264), .A1(n19263), .B0(n19262), .Y(n19286) );
  OAI21XL U4639 ( .A0(n19283), .A1(n19282), .B0(n19281), .Y(n19284) );
  CLKINVX3 U4640 ( .A(n3059), .Y(n8104) );
  OAI21XL U4641 ( .A0(n19237), .A1(n26497), .B0(n14858), .Y(n14938) );
  INVX1 U4642 ( .A(n14939), .Y(n14923) );
  OAI21XL U4643 ( .A0(n14833), .A1(n26504), .B0(n14847), .Y(n14926) );
  OAI21XL U4644 ( .A0(n19237), .A1(n26500), .B0(n14835), .Y(n14946) );
  OAI21XL U4645 ( .A0(n19237), .A1(n25981), .B0(n14857), .Y(n14939) );
  OAI21XL U4646 ( .A0(n19237), .A1(n26507), .B0(n19105), .Y(n19322) );
  INVX1 U4647 ( .A(n19323), .Y(n19278) );
  OAI21XL U4648 ( .A0(n3063), .A1(n26509), .B0(n19214), .Y(n19325) );
  OAI21XL U4649 ( .A0(n19237), .A1(n25957), .B0(n19106), .Y(n19323) );
  OAI21X2 U4650 ( .A0(n3705), .A1(n3704), .B0(n3703), .Y(n16840) );
  INVX4 U4651 ( .A(n7008), .Y(n7364) );
  BUFX4 U4652 ( .A(M0_b_10_), .Y(n25880) );
  OAI21XL U4653 ( .A0(n6274), .A1(n26216), .B0(n6269), .Y(M0_b_4_) );
  OAI21XL U4654 ( .A0(n7422), .A1(n20951), .B0(n3568), .Y(n10729) );
  NOR2X1 U4655 ( .A(n10732), .B(n10734), .Y(n7422) );
  ADDFX2 U4656 ( .A(n16472), .B(n16471), .CI(n16470), .CO(n16464), .S(n16550)
         );
  OAI22X1 U4657 ( .A0(n16962), .A1(n16403), .B0(n16402), .B1(n16960), .Y(
        n16471) );
  INVX8 U4658 ( .A(n2973), .Y(n2974) );
  OAI2BB1X1 U4659 ( .A0N(n17719), .A1N(n3763), .B0(n3762), .Y(n17705) );
  OAI22X1 U4660 ( .A0(n17861), .A1(n17713), .B0(n18141), .B1(n17658), .Y(
        n17719) );
  XNOR2X1 U4661 ( .A(n17965), .B(n3856), .Y(n17997) );
  OAI2BB1X1 U4662 ( .A0N(n17965), .A1N(n3854), .B0(n3853), .Y(n17972) );
  OAI22X1 U4663 ( .A0(n18522), .A1(n17968), .B0(n3195), .B1(n17935), .Y(n17965) );
  OAI22X1 U4664 ( .A0(n16942), .A1(n16516), .B0(n16688), .B1(n16496), .Y(
        n16515) );
  OAI22X1 U4665 ( .A0(n12152), .A1(n11796), .B0(n3185), .B1(n11795), .Y(n11832) );
  OAI2BB2X1 U4666 ( .B0(n3018), .B1(n3685), .A0N(n16113), .A1N(n3684), .Y(
        n16098) );
  OAI22X1 U4667 ( .A0(n16701), .A1(n16107), .B0(n16699), .B1(n16051), .Y(
        n16113) );
  OAI2BB1X1 U4668 ( .A0N(n11845), .A1N(n4421), .B0(n4419), .Y(n12444) );
  OAI22X1 U4669 ( .A0(n12598), .A1(n11850), .B0(n12342), .B1(n11831), .Y(
        n11845) );
  INVXL U4670 ( .A(n10298), .Y(n2975) );
  INVXL U4671 ( .A(n2975), .Y(n2976) );
  ADDFX2 U4672 ( .A(n16796), .B(n16795), .CI(n16794), .CO(n16791), .S(n16829)
         );
  CMPR22X1 U4673 ( .A(n16071), .B(n16070), .CO(n16100), .S(n16795) );
  CMPR22X1 U4674 ( .A(n16355), .B(n16354), .CO(n16391), .S(n16387) );
  OAI22X1 U4675 ( .A0(n17060), .A1(n17038), .B0(n17061), .B1(n16334), .Y(
        n16354) );
  OAI21X1 U4676 ( .A0(n25767), .A1(n26288), .B0(n15943), .Y(M5_a_0_) );
  INVX8 U4677 ( .A(n11479), .Y(n25767) );
  XOR2X1 U4678 ( .A(n12803), .B(n11691), .Y(n3728) );
  INVX1 U4679 ( .A(n2980), .Y(n11691) );
  XNOR2X2 U4680 ( .A(M3_a_10_), .B(M3_a_9_), .Y(n12523) );
  CLKINVX3 U4681 ( .A(M3_a_9_), .Y(n12225) );
  INVX8 U4682 ( .A(n2977), .Y(n2978) );
  CLKINVX3 U4683 ( .A(M3_mult_x_15_a_1_), .Y(n2979) );
  INVX8 U4684 ( .A(n2979), .Y(n2980) );
  NAND2X1 U4685 ( .A(n3389), .B(n3840), .Y(M3_mult_x_15_a_1_) );
  INVXL U4686 ( .A(n24288), .Y(n2981) );
  INVXL U4687 ( .A(n2981), .Y(n2982) );
  CLKINVX3 U4688 ( .A(n2981), .Y(n2983) );
  CLKINVX3 U4689 ( .A(n2981), .Y(n2984) );
  XNOR2XL U4690 ( .A(M2_mult_x_15_a_1_), .B(n9892), .Y(n9902) );
  XNOR2XL U4691 ( .A(n9904), .B(n9892), .Y(n9914) );
  XNOR2XL U4692 ( .A(n21054), .B(n25882), .Y(n6605) );
  XNOR2XL U4693 ( .A(n13049), .B(n13844), .Y(n13093) );
  XNOR2XL U4694 ( .A(n4808), .B(n9960), .Y(n9653) );
  XNOR2XL U4695 ( .A(M2_mult_x_15_a_1_), .B(n10312), .Y(n9844) );
  XNOR2XL U4696 ( .A(M0_b_2_), .B(n3209), .Y(n6616) );
  XNOR2XL U4697 ( .A(n12282), .B(n3110), .Y(n12281) );
  XNOR2XL U4698 ( .A(n25865), .B(n13844), .Y(n13058) );
  XNOR2XL U4699 ( .A(n9904), .B(n10311), .Y(n9815) );
  XNOR2XL U4700 ( .A(n9904), .B(n10341), .Y(n9754) );
  XNOR2XL U4701 ( .A(n25866), .B(n25881), .Y(n6481) );
  XNOR2XL U4702 ( .A(M0_b_2_), .B(n25867), .Y(n6612) );
  XNOR2XL U4703 ( .A(n25867), .B(n7165), .Y(n6479) );
  XNOR2XL U4704 ( .A(n12282), .B(n12271), .Y(n12294) );
  XNOR2XL U4705 ( .A(n3206), .B(M3_mult_x_15_b_3_), .Y(n18149) );
  XNOR2XL U4706 ( .A(M5_mult_x_15_n1), .B(n12279), .Y(n16637) );
  XOR2XL U4707 ( .A(M5_mult_x_15_n1), .B(n3190), .Y(n3792) );
  XNOR2XL U4708 ( .A(n14117), .B(n25860), .Y(n13286) );
  OAI22X1 U4709 ( .A0(n13160), .A1(n13971), .B0(n13172), .B1(n13972), .Y(
        n13166) );
  XNOR2XL U4710 ( .A(n14118), .B(n13844), .Y(n13277) );
  AND2X1 U4711 ( .A(n9937), .B(n9936), .Y(n9938) );
  XNOR2XL U4712 ( .A(n23220), .B(n6944), .Y(n6539) );
  XNOR2XL U4713 ( .A(n4789), .B(n25882), .Y(n6431) );
  XNOR2XL U4714 ( .A(n10494), .B(n9960), .Y(n9599) );
  XOR2XL U4715 ( .A(M3_mult_x_15_b_1_), .B(n3189), .Y(n6096) );
  XNOR2XL U4716 ( .A(n16614), .B(n12279), .Y(n16584) );
  XNOR2XL U4717 ( .A(n16289), .B(n12271), .Y(n16577) );
  XOR2XL U4718 ( .A(n3047), .B(n16965), .Y(n16702) );
  XNOR2XL U4719 ( .A(n13769), .B(n25862), .Y(n13316) );
  XNOR2XL U4720 ( .A(n14266), .B(n13605), .Y(n13391) );
  AND2X1 U4721 ( .A(n13136), .B(n13135), .Y(n13140) );
  NOR2X1 U4722 ( .A(n7382), .B(n26005), .Y(n3475) );
  AOI21XL U4723 ( .A0(n7389), .A1(y10[13]), .B0(n25151), .Y(n4558) );
  ADDFX2 U4724 ( .A(n9995), .B(n9994), .CI(n9993), .CO(n10030), .S(n9997) );
  XNOR2XL U4725 ( .A(n9722), .B(n5746), .Y(n9748) );
  ADDFX2 U4726 ( .A(n9802), .B(n9801), .CI(n9800), .CO(n9810), .S(n10017) );
  XNOR2XL U4727 ( .A(n25868), .B(n25882), .Y(n6363) );
  XNOR2XL U4728 ( .A(n25868), .B(n25881), .Y(n6303) );
  XNOR2XL U4729 ( .A(n21054), .B(M0_b_18_), .Y(n6284) );
  OAI21XL U4730 ( .A0(n6401), .A1(n6402), .B0(n6400), .Y(n3593) );
  ADDFX2 U4731 ( .A(n6520), .B(n6519), .CI(n6518), .CO(n6508), .S(n6640) );
  ADDFX2 U4732 ( .A(n9644), .B(n9643), .CI(n9642), .CO(n9650), .S(n9682) );
  XNOR2XL U4733 ( .A(n12233), .B(n12271), .Y(n12228) );
  XNOR2XL U4734 ( .A(n12519), .B(M3_mult_x_15_b_1_), .Y(n12163) );
  XOR2XL U4735 ( .A(n3198), .B(n4239), .Y(n4877) );
  XNOR2XL U4736 ( .A(n18503), .B(M3_mult_x_15_b_2_), .Y(n18227) );
  XNOR2XL U4737 ( .A(n18118), .B(M3_mult_x_15_b_3_), .Y(n18236) );
  XNOR2XL U4738 ( .A(n18500), .B(M3_mult_x_15_b_2_), .Y(n18050) );
  XNOR2XL U4739 ( .A(n18150), .B(M3_mult_x_15_b_9_), .Y(n18028) );
  AND2X2 U4740 ( .A(n11505), .B(n4480), .Y(n4479) );
  XNOR2XL U4741 ( .A(n16289), .B(M3_mult_x_15_b_6_), .Y(n16531) );
  XNOR2XL U4742 ( .A(n3047), .B(n12561), .Y(n16469) );
  AND2X1 U4743 ( .A(in_valid_t), .B(w2[73]), .Y(n5730) );
  AND3X1 U4744 ( .A(n10799), .B(n10798), .C(n11207), .Y(n22952) );
  XNOR2XL U4745 ( .A(n13769), .B(n14228), .Y(n13403) );
  XNOR2XL U4746 ( .A(n13863), .B(n25862), .Y(n13367) );
  AND2X1 U4747 ( .A(n9101), .B(n5089), .Y(n3454) );
  NOR2X1 U4748 ( .A(n5806), .B(n4108), .Y(n5805) );
  NAND3X1 U4749 ( .A(n9065), .B(n5345), .C(n5344), .Y(M2_a_6_) );
  XNOR2XL U4750 ( .A(n10324), .B(n10342), .Y(n9433) );
  XNOR2XL U4751 ( .A(n25866), .B(n7646), .Y(n6341) );
  XNOR2XL U4752 ( .A(n25867), .B(n7621), .Y(n6735) );
  ADDFX2 U4753 ( .A(n6436), .B(n6435), .CI(n6434), .CO(n6428), .S(n6695) );
  CLKINVX3 U4754 ( .A(n25871), .Y(n6843) );
  INVX1 U4755 ( .A(n6294), .Y(n6295) );
  XOR2XL U4756 ( .A(n12169), .B(n5509), .Y(n12199) );
  XNOR2XL U4757 ( .A(n3204), .B(n12271), .Y(n12341) );
  AND2X1 U4758 ( .A(n12317), .B(n12316), .Y(n12318) );
  XNOR2XL U4759 ( .A(n12233), .B(M3_mult_x_15_b_9_), .Y(n12106) );
  AOI21XL U4760 ( .A0(n4732), .A1(n21166), .B0(n4896), .Y(n4895) );
  NOR2X1 U4761 ( .A(n25796), .B(n26261), .Y(n3880) );
  XNOR2XL U4762 ( .A(n18453), .B(M3_mult_x_15_b_3_), .Y(n17970) );
  XNOR2XL U4763 ( .A(n18118), .B(M3_mult_x_15_b_9_), .Y(n17975) );
  AOI21XL U4764 ( .A0(n11479), .A1(data[98]), .B0(n3677), .Y(n3676) );
  XNOR2XL U4765 ( .A(n16614), .B(n12561), .Y(n16345) );
  AND2X1 U4766 ( .A(n16660), .B(n16659), .Y(n16664) );
  INVX4 U4767 ( .A(n8592), .Y(n3092) );
  OAI21XL U4768 ( .A0(n25243), .A1(n25903), .B0(n11510), .Y(M1_a_4_) );
  NAND3X1 U4769 ( .A(n3286), .B(n3285), .C(n3284), .Y(n3283) );
  AOI21XL U4770 ( .A0(n21166), .A1(n4049), .B0(n5958), .Y(n4048) );
  XNOR2XL U4771 ( .A(n10324), .B(M2_mult_x_15_n1668), .Y(n10158) );
  XNOR2XL U4772 ( .A(n10339), .B(M2_b_15_), .Y(n9345) );
  CLKINVX2 U4773 ( .A(M2_a_3_), .Y(n9907) );
  XNOR2XL U4774 ( .A(n10494), .B(n10312), .Y(n9216) );
  OAI2BB1X1 U4775 ( .A0N(n4730), .A1N(n11536), .B0(n9045), .Y(n6143) );
  XOR2XL U4776 ( .A(n3119), .B(n22492), .Y(n22511) );
  NAND2X1 U4777 ( .A(n25229), .B(target_temp[16]), .Y(n11533) );
  XNOR2XL U4778 ( .A(n23221), .B(n25875), .Y(n7497) );
  XNOR2XL U4779 ( .A(n10494), .B(n9839), .Y(n9204) );
  XOR2XL U4780 ( .A(n10324), .B(n5377), .Y(n5376) );
  AOI21XL U4781 ( .A0(n7389), .A1(y10[20]), .B0(n25157), .Y(n6256) );
  ADDFX2 U4782 ( .A(n6310), .B(n6309), .CI(n6308), .CO(n6796), .S(n6336) );
  BUFX1 U4783 ( .A(n6859), .Y(n4804) );
  XNOR2XL U4784 ( .A(n23220), .B(n7569), .Y(n6922) );
  XNOR2XL U4785 ( .A(n25867), .B(n7646), .Y(n6836) );
  AND2X1 U4786 ( .A(n6662), .B(n6661), .Y(n6663) );
  XOR2X2 U4787 ( .A(n6928), .B(n3591), .Y(n7040) );
  XNOR2XL U4788 ( .A(n23220), .B(n25877), .Y(n7049) );
  XNOR2XL U4789 ( .A(n25869), .B(n25877), .Y(n7149) );
  XNOR2XL U4790 ( .A(n23219), .B(n25875), .Y(n7587) );
  XOR2XL U4791 ( .A(n5970), .B(M3_a_9_), .Y(n3710) );
  XNOR2XL U4792 ( .A(M3_mult_x_15_a_17_), .B(n3049), .Y(n11745) );
  XNOR2XL U4793 ( .A(n12282), .B(n3021), .Y(n12024) );
  ADDFX2 U4794 ( .A(n12143), .B(n12142), .CI(n12141), .CO(n12140), .S(n12177)
         );
  AOI22X2 U4795 ( .A0(n4875), .A1(data[53]), .B0(w2[21]), .B1(in_valid_t), .Y(
        n4441) );
  XOR2XL U4796 ( .A(n18006), .B(M3_mult_x_15_b_20_), .Y(n4188) );
  XNOR2XL U4797 ( .A(n18468), .B(M3_mult_x_15_b_2_), .Y(n17935) );
  XNOR2XL U4798 ( .A(n25864), .B(n25862), .Y(n14046) );
  XOR2XL U4799 ( .A(n3047), .B(n5718), .Y(n16049) );
  ADDFX2 U4800 ( .A(n16398), .B(n16399), .CI(n16400), .CO(n16407), .S(n16465)
         );
  ADDFX2 U4801 ( .A(n16509), .B(n16508), .CI(n16507), .CO(n16555), .S(n16560)
         );
  XOR2X1 U4802 ( .A(M4_a_6_), .B(M4_a_7_), .Y(n4343) );
  XNOR2XL U4803 ( .A(n14236), .B(n14030), .Y(n13600) );
  XNOR2XL U4804 ( .A(n14235), .B(n14030), .Y(n13676) );
  XNOR2XL U4805 ( .A(n14357), .B(n13693), .Y(n13694) );
  CLKINVX3 U4806 ( .A(M1_b_3_), .Y(n13720) );
  INVX4 U4807 ( .A(n6194), .Y(n3016) );
  INVX1 U4808 ( .A(M5_a_18_), .Y(n4797) );
  ADDFX2 U4809 ( .A(n13436), .B(n13435), .CI(n13434), .CO(n13473), .S(n13440)
         );
  INVX4 U4810 ( .A(M2_U4_U1_or2_inv_0__26_), .Y(n9863) );
  CLKINVX2 U4811 ( .A(n4503), .Y(n13280) );
  XNOR2X1 U4812 ( .A(n9477), .B(n5303), .Y(n9472) );
  XOR2XL U4813 ( .A(n4335), .B(n4334), .Y(n9274) );
  NAND3BX1 U4814 ( .AN(n5505), .B(n9079), .C(n5504), .Y(M2_b_13_) );
  NOR2BX2 U4815 ( .AN(n9046), .B(n6143), .Y(n10388) );
  NOR2X2 U4816 ( .A(n3692), .B(n3691), .Y(n16631) );
  XNOR2XL U4817 ( .A(n17039), .B(n12561), .Y(n16201) );
  XNOR2XL U4818 ( .A(n15968), .B(n3202), .Y(n16288) );
  XNOR2XL U4819 ( .A(n25870), .B(n25876), .Y(n7508) );
  ADDFX2 U4820 ( .A(n6761), .B(n6760), .CI(n6759), .CO(n6765), .S(n6770) );
  XOR2X1 U4821 ( .A(n7059), .B(n6992), .Y(n7071) );
  BUFX3 U4822 ( .A(M0_b_5_), .Y(n7164) );
  XNOR2XL U4823 ( .A(n23220), .B(n25874), .Y(n7219) );
  XOR2XL U4824 ( .A(n6288), .B(M0_a_18_), .Y(n6282) );
  XOR2XL U4825 ( .A(n25884), .B(n3201), .Y(n3965) );
  XNOR2XL U4826 ( .A(n25884), .B(n12560), .Y(n11781) );
  XNOR2XL U4827 ( .A(n12594), .B(M3_mult_x_15_b_19_), .Y(n11926) );
  XNOR2XL U4828 ( .A(n12265), .B(n12803), .Y(n11635) );
  XNOR2XL U4829 ( .A(n12265), .B(n3021), .Y(n11847) );
  XNOR2XL U4830 ( .A(n12732), .B(n12279), .Y(n11814) );
  XNOR2XL U4831 ( .A(n12282), .B(n12803), .Y(n11671) );
  XNOR2XL U4832 ( .A(n12233), .B(n12561), .Y(n12033) );
  OAI21X2 U4833 ( .A0(n25913), .A1(n15942), .B0(n4441), .Y(M3_mult_x_15_n61)
         );
  XNOR2XL U4834 ( .A(n18150), .B(n3021), .Y(n17713) );
  ADDFX2 U4835 ( .A(n18040), .B(n18039), .CI(n18038), .CO(n18032), .S(n18101)
         );
  XNOR2XL U4836 ( .A(n18118), .B(n12561), .Y(n17906) );
  XNOR2XL U4837 ( .A(n18500), .B(n3021), .Y(n17558) );
  XNOR2XL U4838 ( .A(n18468), .B(n3048), .Y(n18520) );
  XNOR2XL U4839 ( .A(n15968), .B(n12561), .Y(n16115) );
  XNOR2XL U4840 ( .A(n3203), .B(n3190), .Y(n16063) );
  XOR2XL U4841 ( .A(n5430), .B(n3211), .Y(n3424) );
  XNOR2XL U4842 ( .A(n3047), .B(M3_mult_x_15_b_21_), .Y(n15997) );
  XNOR2XL U4843 ( .A(n3206), .B(n3048), .Y(n17656) );
  BUFX3 U4844 ( .A(n17861), .Y(n18239) );
  AOI21XL U4845 ( .A0(n14417), .A1(y11[18]), .B0(n4771), .Y(n11540) );
  AOI21XL U4846 ( .A0(n19534), .A1(n19771), .B0(n19770), .Y(n19772) );
  CLKINVX3 U4847 ( .A(n14267), .Y(n25863) );
  XNOR2XL U4848 ( .A(n25885), .B(n10386), .Y(n10300) );
  OAI21XL U4849 ( .A0(n25243), .A1(n25899), .B0(n11526), .Y(M1_a_14_) );
  OAI2BB1X1 U4850 ( .A0N(n4111), .A1N(n16447), .B0(n4110), .Y(n16830) );
  BUFX3 U4851 ( .A(M2_b_17_), .Y(n10514) );
  XOR2XL U4852 ( .A(n16972), .B(n5672), .Y(n5671) );
  ADDFX2 U4853 ( .A(n16283), .B(n16282), .CI(n16281), .CO(n16327), .S(n16276)
         );
  NOR2BX1 U4854 ( .AN(n10054), .B(n3091), .Y(n4324) );
  OAI21XL U4855 ( .A0(n6274), .A1(n25994), .B0(n6272), .Y(M0_b_21_) );
  AND2X1 U4856 ( .A(n6726), .B(n6725), .Y(n6727) );
  CLKINVX2 U4857 ( .A(n7695), .Y(n5122) );
  XNOR2XL U4858 ( .A(n12594), .B(M3_mult_x_15_b_22_), .Y(n12596) );
  XNOR2XL U4859 ( .A(n12716), .B(n12560), .Y(n11916) );
  AOI21XL U4860 ( .A0(n3709), .A1(n3665), .B0(n3664), .Y(n3663) );
  XOR2XL U4861 ( .A(M4_a_12_), .B(M4_a_13_), .Y(n5871) );
  XNOR2XL U4862 ( .A(n12758), .B(n3201), .Y(n12553) );
  BUFX3 U4863 ( .A(n12633), .Y(n12513) );
  XNOR2XL U4864 ( .A(n17607), .B(n4488), .Y(n4492) );
  ADDFX2 U4865 ( .A(n3114), .B(n17728), .CI(n17727), .CO(n17760), .S(n17763)
         );
  XNOR2XL U4866 ( .A(n25883), .B(n3190), .Y(n17833) );
  ADDFX2 U4867 ( .A(n14033), .B(n14032), .CI(n14031), .CO(n14063), .S(n14035)
         );
  XOR2XL U4868 ( .A(n16091), .B(n3697), .Y(n3696) );
  OAI2BB1X1 U4869 ( .A0N(n3424), .A1N(n3179), .B0(n3636), .Y(n3635) );
  OAI21XL U4870 ( .A0(n17546), .A1(n17545), .B0(n3432), .Y(n5924) );
  XOR2XL U4871 ( .A(n17568), .B(n3406), .Y(n3405) );
  NOR2X1 U4872 ( .A(n4089), .B(n4088), .Y(n4171) );
  NOR2X1 U4873 ( .A(n14335), .B(n14484), .Y(n14337) );
  AOI21XL U4874 ( .A0(n19936), .A1(n19952), .B0(n3164), .Y(n19935) );
  AND4X1 U4875 ( .A(n8214), .B(n8213), .C(n8212), .D(n8211), .Y(n8215) );
  CLKINVX3 U4876 ( .A(n15161), .Y(n15313) );
  NOR2X1 U4877 ( .A(n23409), .B(n21455), .Y(n21453) );
  AOI21XL U4878 ( .A0(n6202), .A1(n21828), .B0(n21827), .Y(n21829) );
  OAI21XL U4879 ( .A0(n21854), .A1(n21986), .B0(n21985), .Y(n22004) );
  OAI21XL U4880 ( .A0(n3160), .A1(n8802), .B0(n8801), .Y(n8817) );
  XNOR2XL U4881 ( .A(n5677), .B(n3196), .Y(n16892) );
  XNOR2XL U4882 ( .A(n17039), .B(n3048), .Y(n16870) );
  AOI21XL U4883 ( .A0(n10982), .A1(n11005), .B0(n11018), .Y(n10963) );
  XNOR2XL U4884 ( .A(n17073), .B(n3202), .Y(n17059) );
  AOI21XL U4885 ( .A0(n11372), .A1(n11007), .B0(n11023), .Y(n10998) );
  ADDFX2 U4886 ( .A(n10345), .B(n10344), .CI(n10343), .CO(n10414), .S(n10421)
         );
  INVX4 U4887 ( .A(n6014), .Y(n3022) );
  BUFX3 U4888 ( .A(n11487), .Y(M3_mult_x_15_b_19_) );
  NAND2X1 U4889 ( .A(n9508), .B(n9509), .Y(n4118) );
  ADDFX2 U4890 ( .A(n9532), .B(n9531), .CI(n9530), .CO(n9566), .S(n9529) );
  INVX1 U4891 ( .A(n14555), .Y(n4269) );
  ADDFX2 U4892 ( .A(n14147), .B(n14146), .CI(n14145), .CO(n14187), .S(n14144)
         );
  XOR2X1 U4893 ( .A(n3775), .B(n16827), .Y(n16838) );
  NAND3X2 U4894 ( .A(n5189), .B(n4341), .C(n4340), .Y(n5298) );
  OAI21XL U4895 ( .A0(n16045), .A1(n16046), .B0(n16044), .Y(n4152) );
  OAI21XL U4896 ( .A0(n17307), .A1(n17245), .B0(n17246), .Y(n5638) );
  AND2X1 U4897 ( .A(n19278), .B(n19322), .Y(n19279) );
  AOI21X2 U4898 ( .A0(n3512), .A1(n6721), .B0(n6720), .Y(n3511) );
  ADDFX2 U4899 ( .A(n7083), .B(n7082), .CI(n7081), .CO(n7120), .S(n7241) );
  OAI21XL U4900 ( .A0(n7681), .A1(n7745), .B0(n7680), .Y(n7728) );
  XNOR2XL U4901 ( .A(n12732), .B(n12701), .Y(n12639) );
  XOR2XL U4902 ( .A(n4440), .B(n12542), .Y(n4439) );
  XOR2X2 U4903 ( .A(M3_a_11_), .B(n5044), .Y(n12633) );
  OAI21XL U4904 ( .A0(n3928), .A1(n3927), .B0(n3926), .Y(n11822) );
  XNOR2XL U4905 ( .A(n18638), .B(n3048), .Y(n18461) );
  ADDFX2 U4906 ( .A(n17723), .B(n17722), .CI(n17721), .CO(n18343), .S(n18362)
         );
  XNOR2XL U4907 ( .A(n17091), .B(n5053), .Y(n17093) );
  OAI2BB1X1 U4908 ( .A0N(n3868), .A1N(n17705), .B0(n3866), .Y(n17702) );
  OAI2BB1X1 U4909 ( .A0N(n13808), .A1N(n13807), .B0(n13806), .Y(n13809) );
  AOI21XL U4910 ( .A0(n14645), .A1(n14651), .B0(n14344), .Y(n14345) );
  OAI21XL U4911 ( .A0(n3165), .A1(n19936), .B0(n19935), .Y(n19950) );
  NOR2X1 U4912 ( .A(n20377), .B(n8215), .Y(n8598) );
  AOI21XL U4913 ( .A0(n19831), .A1(n19871), .B0(n19830), .Y(n19910) );
  AOI21XL U4914 ( .A0(n20059), .A1(n19891), .B0(n19890), .Y(n19896) );
  INVX4 U4915 ( .A(n15313), .Y(n3090) );
  INVX1 U4916 ( .A(n23125), .Y(n21455) );
  XNOR2XL U4917 ( .A(n21499), .B(n6189), .Y(n21673) );
  AOI21XL U4918 ( .A0(n8702), .A1(n8742), .B0(n8701), .Y(n8781) );
  ADDFX2 U4919 ( .A(n14262), .B(n14261), .CI(n14260), .CO(n14275), .S(n14269)
         );
  OAI2BB1X1 U4920 ( .A0N(n4096), .A1N(n16973), .B0(n4095), .Y(n16969) );
  ADDFX2 U4921 ( .A(n18565), .B(n18564), .CI(n18563), .CO(n18577), .S(n18569)
         );
  ADDFX2 U4922 ( .A(n10360), .B(n10359), .CI(n10358), .CO(n10378), .S(n10424)
         );
  AOI21XL U4923 ( .A0(n17372), .A1(n17139), .B0(n17138), .Y(n17388) );
  XNOR2XL U4924 ( .A(n16953), .B(n16955), .Y(n5687) );
  NAND2X1 U4925 ( .A(n5004), .B(n5003), .Y(n10474) );
  ADDFX2 U4926 ( .A(n14152), .B(n14151), .CI(n14150), .CO(n14184), .S(n14145)
         );
  NAND2X1 U4927 ( .A(n3340), .B(n16077), .Y(n6116) );
  XOR2X1 U4928 ( .A(n16299), .B(n5332), .Y(n16302) );
  NOR2X2 U4929 ( .A(n10124), .B(n10123), .Y(n10201) );
  AOI21XL U4930 ( .A0(n19948), .A1(n20008), .B0(n19947), .Y(n19998) );
  AOI21XL U4931 ( .A0(n15680), .A1(n15511), .B0(n15510), .Y(n15516) );
  XOR2XL U4932 ( .A(n15759), .B(n15755), .Y(n15761) );
  NAND2X1 U4933 ( .A(n10122), .B(n10121), .Y(n10206) );
  OAI2BB1X1 U4934 ( .A0N(n3921), .A1N(n11974), .B0(n3920), .Y(n12683) );
  XOR2X1 U4935 ( .A(n11873), .B(n5975), .Y(n11871) );
  INVX1 U4936 ( .A(n12819), .Y(n4827) );
  AND2X1 U4937 ( .A(n12428), .B(n12427), .Y(n12429) );
  INVX1 U4938 ( .A(n12561), .Y(n12542) );
  AOI21XL U4939 ( .A0(n18993), .A1(n18997), .B0(n18714), .Y(n18715) );
  AND2X1 U4940 ( .A(n18314), .B(n18313), .Y(n18317) );
  AOI21XL U4941 ( .A0(n16760), .A1(n16761), .B0(n16759), .Y(n5657) );
  INVX4 U4942 ( .A(n4210), .Y(n18624) );
  OAI21XL U4943 ( .A0(n13825), .A1(n13826), .B0(n13824), .Y(n6047) );
  XNOR2XL U4944 ( .A(n8896), .B(n8895), .Y(n20439) );
  OAI21XL U4945 ( .A0(n8653), .A1(n8758), .B0(n8652), .Y(n8783) );
  XOR2XL U4946 ( .A(n20062), .B(n20061), .Y(n20186) );
  CLKINVX3 U4947 ( .A(n21580), .Y(n3095) );
  XNOR2XL U4948 ( .A(n22084), .B(n22083), .Y(n22301) );
  AND2X1 U4949 ( .A(n8148), .B(n8192), .Y(n8149) );
  XOR2XL U4950 ( .A(n8767), .B(n8766), .Y(n20461) );
  XNOR2XL U4951 ( .A(n8753), .B(n8752), .Y(n20458) );
  BUFX8 U4952 ( .A(M3_mult_x_15_b_22_), .Y(n3202) );
  NOR2X1 U4953 ( .A(n14320), .B(n14319), .Y(n14160) );
  ADDFX2 U4954 ( .A(n17054), .B(n17055), .CI(n17053), .CO(n17067), .S(n17062)
         );
  INVX1 U4955 ( .A(n10467), .Y(n3150) );
  ADDFX2 U4956 ( .A(n16899), .B(n16898), .CI(n16897), .CO(n16915), .S(n16900)
         );
  ADDFX2 U4957 ( .A(n17049), .B(n17048), .CI(n17047), .CO(n17050), .S(n17033)
         );
  OAI21X1 U4958 ( .A0(n5077), .A1(n4175), .B0(n3829), .Y(n3828) );
  OAI2BB1X1 U4959 ( .A0N(n5331), .A1N(n16299), .B0(n5330), .Y(n17016) );
  NAND2X1 U4960 ( .A(n10124), .B(n10123), .Y(n10202) );
  OAI21X1 U4961 ( .A0(n5602), .A1(n10735), .B0(n20951), .Y(n3482) );
  XOR2XL U4962 ( .A(n15684), .B(n15683), .Y(n15809) );
  NOR2X1 U4963 ( .A(n12776), .B(n12777), .Y(n12841) );
  AOI21X2 U4964 ( .A0(n3888), .A1(n3889), .B0(n12429), .Y(n3887) );
  ADDFX2 U4965 ( .A(n18443), .B(n18442), .CI(n18441), .CO(n18459), .S(n18513)
         );
  XNOR2XL U4966 ( .A(n18722), .B(n3202), .Y(n18723) );
  OAI21XL U4967 ( .A0(n18692), .A1(n18927), .B0(n18691), .Y(n18693) );
  XNOR2XL U4968 ( .A(n19882), .B(n19881), .Y(n20255) );
  XOR2XL U4969 ( .A(n9000), .B(n8999), .Y(n9006) );
  OAI21XL U4970 ( .A0(n3067), .A1(n9002), .B0(n9001), .Y(n9005) );
  XOR2XL U4971 ( .A(n20043), .B(n20042), .Y(n20195) );
  XOR2XL U4972 ( .A(n20147), .B(n20141), .Y(n20149) );
  OAI21XL U4973 ( .A0(n3030), .A1(n20143), .B0(n20142), .Y(n20148) );
  OAI21XL U4974 ( .A0(n21386), .A1(n21385), .B0(n21384), .Y(n21387) );
  OAI21XL U4975 ( .A0(n14833), .A1(n26503), .B0(n14849), .Y(n14954) );
  XNOR2XL U4976 ( .A(n22056), .B(n22055), .Y(n22254) );
  OR2X2 U4977 ( .A(n21737), .B(n3222), .Y(n21854) );
  INVX4 U4978 ( .A(n11536), .Y(n3103) );
  NAND2X1 U4979 ( .A(n12503), .B(n12502), .Y(n12887) );
  NOR2X1 U4980 ( .A(n17109), .B(n17108), .Y(n17316) );
  INVX1 U4981 ( .A(n14160), .Y(n14526) );
  NOR2X2 U4982 ( .A(n10128), .B(n10129), .Y(n10218) );
  NOR2X1 U4983 ( .A(n14545), .B(n14529), .Y(n14535) );
  NOR2X1 U4984 ( .A(n14326), .B(n14325), .Y(n14545) );
  NAND2X1 U4985 ( .A(n10133), .B(n10132), .Y(n10244) );
  AOI21XL U4986 ( .A0(n10597), .A1(n10601), .B0(n10579), .Y(n10580) );
  AND2X1 U4987 ( .A(n5032), .B(data[60]), .Y(n11571) );
  INVX1 U4988 ( .A(n3310), .Y(n3233) );
  AOI21XL U4989 ( .A0(n19286), .A1(n19285), .B0(n19284), .Y(n19287) );
  AND2X1 U4990 ( .A(n25206), .B(data[62]), .Y(n11553) );
  NAND2X1 U4991 ( .A(n7263), .B(n7262), .Y(n7424) );
  AOI21XL U4992 ( .A0(n7704), .A1(n7703), .B0(n7702), .Y(n7705) );
  AND2X1 U4993 ( .A(n7867), .B(n10726), .Y(n4673) );
  NOR2X2 U4994 ( .A(n12992), .B(n4700), .Y(n3985) );
  NAND2X2 U4995 ( .A(n4035), .B(n4034), .Y(n12865) );
  NAND2X1 U4996 ( .A(n18393), .B(n18392), .Y(n18728) );
  AND2X1 U4997 ( .A(n18955), .B(n18956), .Y(n4639) );
  NAND2X2 U4998 ( .A(n20970), .B(n3737), .Y(n3446) );
  ADDFX2 U4999 ( .A(n18628), .B(n18627), .CI(n18626), .CO(n18629), .S(n18616)
         );
  XOR2XL U5000 ( .A(n19027), .B(n19026), .Y(n18778) );
  INVX1 U5001 ( .A(n20378), .Y(n8179) );
  XNOR2XL U5002 ( .A(n15591), .B(n15590), .Y(n24962) );
  OAI21XL U5003 ( .A0(n8154), .A1(n8153), .B0(n8152), .Y(n8155) );
  OAI21X1 U5004 ( .A0(n14677), .A1(n14590), .B0(n14591), .Y(n14577) );
  AND2X1 U5005 ( .A(n18847), .B(n18848), .Y(n18849) );
  XOR2X1 U5006 ( .A(n10573), .B(n4703), .Y(n20714) );
  NOR2X2 U5007 ( .A(n23736), .B(n23739), .Y(n19098) );
  NOR2X1 U5008 ( .A(n6142), .B(n20646), .Y(n5247) );
  NAND2X1 U5009 ( .A(n16863), .B(n16862), .Y(n17307) );
  OAI21XL U5010 ( .A0(n3041), .A1(n19332), .B0(n19331), .Y(n23209) );
  NOR2X2 U5011 ( .A(n19058), .B(n19077), .Y(n20894) );
  CLKINVX3 U5012 ( .A(n3127), .Y(n3070) );
  AND2X1 U5013 ( .A(n10703), .B(n20944), .Y(n4353) );
  INVX1 U5014 ( .A(n12770), .Y(n4910) );
  CLKINVX3 U5015 ( .A(n22395), .Y(n22343) );
  OAI21XL U5016 ( .A0(n26144), .A1(n21333), .B0(n21332), .Y(n21413) );
  CLKINVX3 U5017 ( .A(n22188), .Y(n22308) );
  INVX1 U5018 ( .A(n3934), .Y(n3338) );
  AOI21XL U5019 ( .A0(n3223), .A1(sigma10[29]), .B0(n14415), .Y(n14707) );
  AND2X1 U5020 ( .A(n17318), .B(n17317), .Y(n4638) );
  XOR2X1 U5021 ( .A(n5139), .B(n4606), .Y(n23495) );
  XOR2X1 U5022 ( .A(n14677), .B(n14593), .Y(n23447) );
  XOR2X1 U5023 ( .A(n4406), .B(n18916), .Y(n23458) );
  NAND2X1 U5024 ( .A(n20709), .B(n20710), .Y(n4245) );
  XOR2XL U5025 ( .A(n11580), .B(n13007), .Y(n11606) );
  AND2X1 U5026 ( .A(n20371), .B(n20372), .Y(n20368) );
  XOR2XL U5027 ( .A(n7446), .B(n6959), .Y(n19076) );
  XOR2XL U5028 ( .A(n7843), .B(n7842), .Y(n7409) );
  AOI21XL U5029 ( .A0(n12835), .A1(n12858), .B0(n12859), .Y(n12860) );
  NAND2X1 U5030 ( .A(n20317), .B(n20315), .Y(n21022) );
  CLKINVX2 U5031 ( .A(n19020), .Y(n23519) );
  AND2X2 U5032 ( .A(n4197), .B(n5439), .Y(n3837) );
  XOR2XL U5033 ( .A(n14433), .B(n14707), .Y(n14458) );
  INVX1 U5034 ( .A(n20838), .Y(n24789) );
  INVX1 U5035 ( .A(n24813), .Y(n24760) );
  OAI21XL U5036 ( .A0(n23957), .A1(n23956), .B0(n23955), .Y(n23961) );
  AOI21XL U5037 ( .A0(n14904), .A1(n14903), .B0(n14902), .Y(n14905) );
  INVX4 U5038 ( .A(n11483), .Y(n5480) );
  XOR2X2 U5039 ( .A(n3795), .B(n4638), .Y(n17425) );
  INVX1 U5040 ( .A(n17435), .Y(n20355) );
  XOR2X1 U5041 ( .A(n3807), .B(n4630), .Y(n17467) );
  AND2X1 U5042 ( .A(n13023), .B(n19042), .Y(n23078) );
  XNOR2XL U5043 ( .A(n24575), .B(n24574), .Y(n24576) );
  NAND2X1 U5044 ( .A(n15793), .B(n15786), .Y(n15818) );
  XOR2XL U5045 ( .A(n20881), .B(n20880), .Y(n23580) );
  NAND2X1 U5046 ( .A(n7871), .B(n4689), .Y(n5569) );
  XNOR2XL U5047 ( .A(n20916), .B(n20915), .Y(n20917) );
  XOR2XL U5048 ( .A(n20851), .B(n20850), .Y(n20852) );
  INVX1 U5049 ( .A(n23760), .Y(n23761) );
  XNOR2XL U5050 ( .A(n24789), .B(n23581), .Y(n23582) );
  XNOR2XL U5051 ( .A(n24760), .B(n24596), .Y(n24597) );
  XOR2XL U5052 ( .A(n20263), .B(n24688), .Y(n20264) );
  XOR2XL U5053 ( .A(n24954), .B(n25353), .Y(n24955) );
  XOR2XL U5054 ( .A(n25288), .B(n25287), .Y(n25289) );
  AOI21X2 U5055 ( .A0(n23963), .A1(n15794), .B0(n4451), .Y(n24428) );
  INVX1 U5056 ( .A(in_valid_w1), .Y(n21110) );
  XNOR2XL U5057 ( .A(n23295), .B(n23294), .Y(n23296) );
  XOR2XL U5058 ( .A(n23309), .B(n23308), .Y(n23310) );
  BUFX3 U5059 ( .A(n23255), .Y(n23256) );
  OAI21XL U5060 ( .A0(n19237), .A1(n25246), .B0(n8217), .Y(n23176) );
  XOR2XL U5061 ( .A(n23712), .B(n23711), .Y(n23881) );
  XOR2XL U5062 ( .A(n21036), .B(n23572), .Y(n24183) );
  XOR2X1 U5063 ( .A(n20741), .B(n20740), .Y(n20936) );
  XOR2X1 U5064 ( .A(n23490), .B(n23736), .Y(n23944) );
  XOR2XL U5065 ( .A(n3456), .B(n20893), .Y(n23619) );
  NAND2X1 U5066 ( .A(n23723), .B(n3128), .Y(n5482) );
  AOI22X1 U5067 ( .A0(n3455), .A1(n20872), .B0(n23893), .B1(n3139), .Y(n23593)
         );
  XOR2XL U5068 ( .A(n22466), .B(n22465), .Y(n23041) );
  XNOR2XL U5069 ( .A(n24503), .B(n24483), .Y(n24484) );
  XNOR2XL U5070 ( .A(n24557), .B(n24556), .Y(n24558) );
  XOR2XL U5071 ( .A(n24778), .B(n24777), .Y(n24779) );
  XOR2XL U5072 ( .A(n24978), .B(n25281), .Y(n24979) );
  XOR2XL U5073 ( .A(n20854), .B(n20866), .Y(n20899) );
  NOR2X1 U5074 ( .A(n7871), .B(n7870), .Y(n23868) );
  XOR2XL U5075 ( .A(n24262), .B(n20695), .Y(n24263) );
  XOR2X2 U5076 ( .A(n4523), .B(n4685), .Y(n5899) );
  NAND3BX1 U5077 ( .AN(n4093), .B(n4094), .C(n25767), .Y(n25757) );
  NAND2X1 U5078 ( .A(n22228), .B(n22217), .Y(n23235) );
  AOI22X1 U5079 ( .A0(n23881), .A1(n3081), .B0(n5340), .B1(n4267), .Y(n24847)
         );
  AOI21XL U5080 ( .A0(n23769), .A1(n3066), .B0(n4843), .Y(n23931) );
  AOI21XL U5081 ( .A0(n23758), .A1(n3066), .B0(n4872), .Y(n20827) );
  AOI21XL U5082 ( .A0(n24526), .A1(n3123), .B0(n23474), .Y(n23475) );
  AOI21XL U5083 ( .A0(n3602), .A1(n3065), .B0(n20631), .Y(n20632) );
  OAI21XL U5084 ( .A0(n25556), .A1(n20748), .B0(n24553), .Y(n24554) );
  OAI21XL U5085 ( .A0(n24352), .A1(n3024), .B0(n24345), .Y(n24346) );
  OAI2BB1X2 U5086 ( .A0N(n23534), .A1N(n19075), .B0(n5482), .Y(n19089) );
  INVX1 U5087 ( .A(n23593), .Y(n24677) );
  OAI21XL U5088 ( .A0(n24439), .A1(n24393), .B0(n24392), .Y(n24459) );
  OAI21XL U5089 ( .A0(n24439), .A1(n24075), .B0(n24074), .Y(n24414) );
  NAND2X1 U5090 ( .A(n3489), .B(n3488), .Y(n23769) );
  AND2X1 U5091 ( .A(n24211), .B(n4950), .Y(n24214) );
  XOR2X1 U5092 ( .A(n5900), .B(n5899), .Y(n24244) );
  NOR2X2 U5093 ( .A(n26140), .B(cs[1]), .Y(n23970) );
  OAI2BB1X1 U5094 ( .A0N(n17436), .A1N(n3136), .B0(n5721), .Y(mul5_out[13]) );
  OAI2BB1X1 U5095 ( .A0N(n25807), .A1N(n24673), .B0(n3530), .Y(n2592) );
  AOI21XL U5096 ( .A0(n24677), .A1(n3060), .B0(n24676), .Y(n2416) );
  AOI21XL U5097 ( .A0(n23579), .A1(n3060), .B0(n23578), .Y(n2410) );
  AOI21XL U5098 ( .A0(n24606), .A1(n3060), .B0(n24605), .Y(n2409) );
  AOI21XL U5099 ( .A0(n5408), .A1(n20353), .B0(n21026), .Y(n2268) );
  AOI21XL U5100 ( .A0(n4893), .A1(n25767), .B0(n25766), .Y(n2286) );
  OAI21XL U5101 ( .A0(mul5_out[0]), .A1(n4772), .B0(n24265), .Y(n2296) );
  CLKINVX2 U5102 ( .A(n4581), .Y(n3065) );
  INVX4 U5103 ( .A(in_valid_d), .Y(n4580) );
  INVX4 U5104 ( .A(n3103), .Y(n25233) );
  CLKINVX2 U5105 ( .A(in_valid_d), .Y(n4585) );
  AND2X1 U5106 ( .A(n11479), .B(data[105]), .Y(n2987) );
  AND2X1 U5107 ( .A(n23556), .B(n23548), .Y(n2988) );
  OR2X2 U5108 ( .A(n24188), .B(n4586), .Y(n2990) );
  XOR2X2 U5109 ( .A(n3415), .B(n12913), .Y(n13029) );
  AND2X2 U5110 ( .A(n23513), .B(n23515), .Y(n2991) );
  CLKINVX2 U5111 ( .A(n3021), .Y(n3043) );
  XNOR2XL U5112 ( .A(n3047), .B(n4206), .Y(n2992) );
  BUFX1 U5113 ( .A(n5437), .Y(n4197) );
  CLKINVX3 U5114 ( .A(n5437), .Y(n4198) );
  INVX4 U5115 ( .A(n4002), .Y(n12265) );
  XOR2X2 U5116 ( .A(n4379), .B(n12832), .Y(n13037) );
  INVX4 U5117 ( .A(n18658), .Y(n25883) );
  NAND2X4 U5118 ( .A(n14356), .B(n13609), .Y(n2993) );
  AND2X2 U5119 ( .A(n9071), .B(n3559), .Y(n2994) );
  INVX1 U5120 ( .A(n21849), .Y(n21859) );
  AND2X2 U5121 ( .A(n3222), .B(n21737), .Y(n21849) );
  INVX1 U5122 ( .A(n6288), .Y(n7644) );
  INVX4 U5123 ( .A(n10388), .Y(M2_mult_x_15_n43) );
  INVX1 U5124 ( .A(n23548), .Y(n23558) );
  CLKINVX3 U5125 ( .A(n25542), .Y(n3228) );
  CLKBUFX8 U5126 ( .A(n25567), .Y(n3061) );
  OR3XL U5127 ( .A(n9043), .B(n25696), .C(n2972), .Y(n23764) );
  CLKINVX2 U5128 ( .A(n13051), .Y(n14029) );
  OR2X2 U5129 ( .A(n15941), .B(n6203), .Y(n2995) );
  XOR2X2 U5130 ( .A(n19357), .B(n19356), .Y(n2996) );
  INVX4 U5131 ( .A(n3166), .Y(n3035) );
  NAND2X4 U5132 ( .A(n13044), .B(n13899), .Y(n2997) );
  CLKBUFX8 U5133 ( .A(M4_mult_x_15_n1680), .Y(n16884) );
  INVX1 U5134 ( .A(n14120), .Y(n13203) );
  NOR2X2 U5135 ( .A(n25567), .B(n3026), .Y(n21113) );
  NAND2X1 U5136 ( .A(n10329), .B(n5078), .Y(n10548) );
  BUFX1 U5137 ( .A(n11479), .Y(n5015) );
  CLKINVX2 U5138 ( .A(n25813), .Y(n4772) );
  INVX4 U5139 ( .A(n12731), .Y(n12732) );
  CLKINVX2 U5140 ( .A(n4945), .Y(n12731) );
  INVX12 U5141 ( .A(n25584), .Y(n3216) );
  CLKINVX3 U5142 ( .A(n25541), .Y(n25584) );
  AND2X1 U5143 ( .A(cs[0]), .B(cs[1]), .Y(n4631) );
  CLKINVX3 U5144 ( .A(n4631), .Y(n21329) );
  AND2X2 U5145 ( .A(n6015), .B(n6017), .Y(n6014) );
  CLKINVX2 U5146 ( .A(M4_a_7_), .Y(n18106) );
  AOI21XL U5147 ( .A0(n8936), .A1(n8935), .B0(n8934), .Y(n9003) );
  CLKINVX3 U5148 ( .A(n3079), .Y(n3130) );
  INVX1 U5149 ( .A(n3599), .Y(n6293) );
  XOR2X1 U5150 ( .A(n5682), .B(n4692), .Y(n17469) );
  CLKINVX3 U5151 ( .A(n15808), .Y(n3125) );
  INVX4 U5152 ( .A(n3709), .Y(n12598) );
  AND2X2 U5153 ( .A(n3710), .B(n12342), .Y(n3709) );
  ADDFX2 U5154 ( .A(n9291), .B(n9290), .CI(n9289), .CO(n9368), .S(n9292) );
  XNOR2X2 U5155 ( .A(n15970), .B(M5_a_2_), .Y(n5835) );
  NAND2X1 U5156 ( .A(n11624), .B(n12284), .Y(n12025) );
  OR2X2 U5157 ( .A(n16727), .B(n16726), .Y(n2998) );
  INVX4 U5158 ( .A(M3_U3_U1_or2_inv_0__18_), .Y(n12519) );
  XNOR2X4 U5159 ( .A(n3884), .B(n4612), .Y(n2999) );
  NOR2X1 U5160 ( .A(n12774), .B(n12775), .Y(n12848) );
  OAI21X2 U5161 ( .A0(n12981), .A1(n3844), .B0(n12982), .Y(n12835) );
  INVX1 U5162 ( .A(n12835), .Y(n12851) );
  OR2X2 U5163 ( .A(n18684), .B(n18683), .Y(n3000) );
  XNOR2X1 U5164 ( .A(n20357), .B(n17466), .Y(n3001) );
  AND2X2 U5165 ( .A(n3933), .B(n17435), .Y(n3002) );
  NOR2X2 U5166 ( .A(n12506), .B(n12505), .Y(n12906) );
  ADDFX2 U5167 ( .A(n13931), .B(n13930), .CI(n13929), .CO(n13979), .S(n13936)
         );
  NOR2X1 U5168 ( .A(n13594), .B(n5258), .Y(n14398) );
  BUFX1 U5169 ( .A(n6298), .Y(n5596) );
  CLKINVX3 U5170 ( .A(n5596), .Y(n7460) );
  INVX4 U5171 ( .A(n18428), .Y(n18500) );
  NOR2X2 U5172 ( .A(n3783), .B(n3782), .Y(n16873) );
  INVX1 U5173 ( .A(n12891), .Y(n12919) );
  AND2X2 U5174 ( .A(n4501), .B(n4500), .Y(n3004) );
  AND2X2 U5175 ( .A(n4501), .B(n4499), .Y(n3005) );
  AND3X4 U5176 ( .A(n23551), .B(n3354), .C(n4222), .Y(n3006) );
  AND2X2 U5177 ( .A(n4408), .B(n18791), .Y(n3007) );
  INVX4 U5178 ( .A(n4227), .Y(n17512) );
  XOR2X1 U5179 ( .A(n5470), .B(n18658), .Y(n4227) );
  OAI21X1 U5180 ( .A0(n18890), .A1(n18899), .B0(n18891), .Y(n18867) );
  NOR2X2 U5181 ( .A(n3625), .B(n3624), .Y(n4796) );
  INVX1 U5182 ( .A(n17431), .Y(n5719) );
  XOR2X2 U5183 ( .A(n4130), .B(n17333), .Y(n17431) );
  NAND2X1 U5184 ( .A(n10118), .B(n10117), .Y(n10280) );
  XNOR2X2 U5185 ( .A(n10065), .B(n4468), .Y(n3008) );
  OAI21XL U5186 ( .A0(n5223), .A1(n5222), .B0(n5221), .Y(n10428) );
  CLKINVX2 U5187 ( .A(n19952), .Y(n3215) );
  AND2X2 U5188 ( .A(n3852), .B(n3085), .Y(n3009) );
  INVX1 U5189 ( .A(n3627), .Y(n5848) );
  INVX1 U5190 ( .A(n17427), .Y(n3627) );
  AND3X1 U5191 ( .A(n17443), .B(n20744), .C(n17450), .Y(n3010) );
  AND2X2 U5192 ( .A(n20808), .B(n4306), .Y(n3011) );
  NOR2X2 U5193 ( .A(n10141), .B(n10140), .Y(n10195) );
  INVX4 U5194 ( .A(n3071), .Y(n3031) );
  XOR2X1 U5195 ( .A(n10196), .B(n4640), .Y(n23533) );
  CLKINVX2 U5196 ( .A(n23533), .Y(n3817) );
  OR2X2 U5197 ( .A(n7815), .B(n7821), .Y(n3012) );
  XOR2X2 U5198 ( .A(n3552), .B(n4680), .Y(n20757) );
  AND2X2 U5199 ( .A(n20869), .B(n20853), .Y(n3013) );
  INVX1 U5200 ( .A(n20284), .Y(n20366) );
  NOR2X1 U5201 ( .A(n20760), .B(n20284), .Y(n3537) );
  INVX4 U5202 ( .A(n3101), .Y(n15190) );
  AOI21XL U5203 ( .A0(n19072), .A1(n24525), .B0(n24471), .Y(n2395) );
  INVX1 U5204 ( .A(n24817), .Y(n25435) );
  AOI22XL U5205 ( .A0(n24692), .A1(n24807), .B0(n24908), .B1(n24764), .Y(
        n24765) );
  AOI22XL U5206 ( .A0(n24692), .A1(n24951), .B0(n24908), .B1(n24863), .Y(
        n24864) );
  AOI22XL U5207 ( .A0(n24692), .A1(n24950), .B0(n24908), .B1(n24907), .Y(
        n24909) );
  AOI22XL U5208 ( .A0(n24692), .A1(n24956), .B0(n24908), .B1(n24955), .Y(
        n24957) );
  AOI22X1 U5209 ( .A0(n3029), .A1(n24469), .B0(n25290), .B1(n24468), .Y(n25625) );
  AOI22XL U5210 ( .A0(n24692), .A1(n24808), .B0(n24908), .B1(n24730), .Y(
        n24731) );
  AOI21XL U5211 ( .A0(n3550), .A1(n24525), .B0(n25031), .Y(n2434) );
  AOI22XL U5212 ( .A0(n24570), .A1(n24692), .B0(n24908), .B1(n24551), .Y(
        n24552) );
  AOI21X1 U5213 ( .A0(n6161), .A1(n3602), .B0(n23842), .Y(n2432) );
  INVX1 U5214 ( .A(n24675), .Y(n25486) );
  AOI222XL U5215 ( .A0(n25745), .A1(n25744), .B0(n25743), .B1(y20[0]), .C0(
        n25742), .C1(n20890), .Y(n2360) );
  AOI222XL U5216 ( .A0(n23769), .A1(n25744), .B0(n25743), .B1(y20[8]), .C0(
        n25535), .C1(n20890), .Y(n2368) );
  AOI222XL U5217 ( .A0(n24514), .A1(n25744), .B0(n25743), .B1(y20[3]), .C0(
        n25597), .C1(n20890), .Y(n2363) );
  NAND2X2 U5218 ( .A(n20172), .B(n20171), .Y(n20194) );
  XOR2XL U5219 ( .A(n24791), .B(n4778), .Y(n24792) );
  INVX1 U5220 ( .A(n24687), .Y(n24726) );
  INVX1 U5221 ( .A(n24980), .Y(n25281) );
  NAND2X4 U5222 ( .A(n20382), .B(n20381), .Y(n20425) );
  NAND2X1 U5223 ( .A(n24541), .B(n24518), .Y(n24583) );
  NOR2X1 U5224 ( .A(n20493), .B(n24784), .Y(n20516) );
  XOR2X1 U5225 ( .A(n23372), .B(n23371), .Y(n23373) );
  OR2X2 U5226 ( .A(n20243), .B(n20066), .Y(n24835) );
  AOI2BB2X1 U5227 ( .B0(n24301), .B1(n20129), .A0N(n20129), .A1N(n24301), .Y(
        n24299) );
  AOI2BB2XL U5228 ( .B0(n24018), .B1(n15739), .A0N(n15739), .A1N(n24018), .Y(
        n24019) );
  NOR2X1 U5229 ( .A(n24877), .B(n15638), .Y(n24502) );
  INVX1 U5230 ( .A(n20380), .Y(n20381) );
  NAND2X1 U5231 ( .A(n23625), .B(n20898), .Y(n24561) );
  NOR2X1 U5232 ( .A(n20519), .B(n8997), .Y(n24566) );
  NOR2X1 U5233 ( .A(n20602), .B(n8997), .Y(n20898) );
  NOR2X1 U5234 ( .A(n20590), .B(n8997), .Y(n23625) );
  OAI22X1 U5235 ( .A0(n3072), .A1(n20211), .B0(n20148), .B1(n3032), .Y(n20181)
         );
  NOR2X1 U5236 ( .A(n20574), .B(n8997), .Y(n20913) );
  XOR2X1 U5237 ( .A(n23280), .B(n23279), .Y(n23281) );
  ADDFHX1 U5238 ( .A(n24296), .B(n3074), .CI(n20122), .CO(n20121), .S(n24294)
         );
  NOR2X1 U5239 ( .A(n20552), .B(n8997), .Y(n23773) );
  NAND2X1 U5240 ( .A(n3030), .B(n20156), .Y(n20139) );
  NAND2X1 U5241 ( .A(n3030), .B(n20149), .Y(n20142) );
  NAND2X1 U5242 ( .A(n23318), .B(n23322), .Y(n23344) );
  NOR2X1 U5243 ( .A(n20533), .B(n20532), .Y(n20591) );
  NOR2X1 U5244 ( .A(n15764), .B(n23956), .Y(n15765) );
  OAI22X1 U5245 ( .A0(n9012), .A1(n3031), .B0(n9006), .B1(n3071), .Y(n20512)
         );
  AOI2BB2XL U5246 ( .B0(n20505), .B1(n3068), .A0N(n20504), .A1N(n3068), .Y(
        n20556) );
  NOR2X1 U5247 ( .A(n22446), .B(n23113), .Y(n23277) );
  INVX2 U5248 ( .A(n20125), .Y(n24986) );
  AOI2BB2X1 U5249 ( .B0(n23397), .B1(n22173), .A0N(n22173), .A1N(n23397), .Y(
        n23396) );
  NAND2BXL U5250 ( .AN(n23942), .B(n4829), .Y(n4828) );
  NOR2X1 U5251 ( .A(n22279), .B(n22278), .Y(n22342) );
  NOR2X1 U5252 ( .A(n3126), .B(n22306), .Y(n22310) );
  AOI21X1 U5253 ( .A0(n24548), .A1(n3123), .B0(n23890), .Y(n23891) );
  INVX4 U5254 ( .A(n20138), .Y(n3072) );
  NAND2BXL U5255 ( .AN(n23889), .B(n23888), .Y(n23890) );
  NAND2X1 U5256 ( .A(n23409), .B(n22188), .Y(n22179) );
  NAND2X1 U5257 ( .A(n4240), .B(n24180), .Y(n24181) );
  AOI22XL U5258 ( .A0(n24397), .A1(n25807), .B0(n2983), .B1(temp2[28]), .Y(
        n24398) );
  NAND3X1 U5259 ( .A(n23570), .B(n23571), .C(n6048), .Y(n2549) );
  NAND2XL U5260 ( .A(n24535), .B(in_valid_d), .Y(n6048) );
  NAND3X1 U5261 ( .A(n3128), .B(n20950), .C(n3050), .Y(n3315) );
  INVXL U5262 ( .A(n24277), .Y(n25168) );
  NAND2XL U5263 ( .A(n5821), .B(n24207), .Y(n24208) );
  AOI21X1 U5264 ( .A0(n24555), .A1(n3066), .B0(n4716), .Y(n4992) );
  OAI21X1 U5265 ( .A0(n4380), .A1(n4772), .B0(n25751), .Y(n25752) );
  OAI21X2 U5266 ( .A0(n5914), .A1(n20786), .B0(n4173), .Y(n20659) );
  AOI22X1 U5267 ( .A0(n4215), .A1(n5017), .B0(n25379), .B1(n4220), .Y(n4380)
         );
  NAND2XL U5268 ( .A(n24199), .B(n5269), .Y(n5268) );
  OAI2BB1XL U5269 ( .A0N(n24117), .A1N(n25527), .B0(n24152), .Y(n24153) );
  NAND2BX1 U5270 ( .AN(n24595), .B(n3065), .Y(n3459) );
  NOR2X1 U5271 ( .A(n20771), .B(n20769), .Y(n20765) );
  NAND2XL U5272 ( .A(n25378), .B(n3080), .Y(n3408) );
  AOI22XL U5273 ( .A0(n5017), .A1(n25638), .B0(n2983), .B1(temp2[22]), .Y(
        n23555) );
  INVX1 U5274 ( .A(n5017), .Y(n25758) );
  INVXL U5275 ( .A(n24244), .Y(n24233) );
  OAI21XL U5276 ( .A0(mul5_out[19]), .A1(n4772), .B0(n4854), .Y(n2334) );
  OAI21XL U5277 ( .A0(n25757), .A1(n24255), .B0(n24054), .Y(n24055) );
  OAI21XL U5278 ( .A0(mul5_out[18]), .A1(n4772), .B0(n4853), .Y(n2332) );
  CLKINVX3 U5279 ( .A(n25757), .Y(n3080) );
  NOR2X1 U5280 ( .A(n25328), .B(n25330), .Y(n25297) );
  NOR2BX1 U5281 ( .AN(n24220), .B(n25328), .Y(n24223) );
  OAI21XL U5282 ( .A0(mul5_out[9]), .A1(n3111), .B0(n24159), .Y(n2314) );
  OAI21XL U5283 ( .A0(mul5_out[12]), .A1(n5434), .B0(n24182), .Y(n2320) );
  OAI21XL U5284 ( .A0(mul5_out[16]), .A1(n4772), .B0(n24219), .Y(n2328) );
  OAI21XL U5285 ( .A0(mul5_out[8]), .A1(n4772), .B0(n20339), .Y(n2312) );
  OAI21XL U5286 ( .A0(mul5_out[7]), .A1(n3111), .B0(n4849), .Y(n2310) );
  OAI21XL U5287 ( .A0(mul5_out[5]), .A1(n3111), .B0(n24134), .Y(n2306) );
  AOI2BB1XL U5288 ( .A0N(n22148), .A1N(n22285), .B0(n22282), .Y(n22149) );
  NAND2XL U5289 ( .A(n3975), .B(n3974), .Y(n3973) );
  INVXL U5290 ( .A(n15782), .Y(n15783) );
  INVX1 U5291 ( .A(n24962), .Y(n3133) );
  AOI2BB1XL U5292 ( .A0N(n22147), .A1N(n22287), .B0(n22286), .Y(n22148) );
  NAND2X1 U5293 ( .A(n20942), .B(n5336), .Y(n5949) );
  NAND2X1 U5294 ( .A(n20942), .B(n3136), .Y(n5851) );
  NAND2XL U5295 ( .A(n23565), .B(n20697), .Y(n5425) );
  INVX1 U5296 ( .A(n24783), .Y(n25735) );
  NOR2XL U5297 ( .A(n25331), .B(n25330), .Y(n25334) );
  NAND2X1 U5298 ( .A(n23744), .B(n20974), .Y(n20976) );
  NOR2X2 U5299 ( .A(n3140), .B(n5033), .Y(n4524) );
  AOI2BB1XL U5300 ( .A0N(n20083), .A1N(n20204), .B0(n20203), .Y(n20084) );
  NOR2XL U5301 ( .A(n23732), .B(n3859), .Y(n3858) );
  AND2X1 U5302 ( .A(n24252), .B(n24253), .Y(n25637) );
  INVX4 U5303 ( .A(n23734), .Y(n3014) );
  AOI21XL U5304 ( .A0(n25220), .A1(n25108), .B0(n25219), .Y(n25109) );
  NAND2XL U5305 ( .A(n23732), .B(n4222), .Y(n4216) );
  NAND2X1 U5306 ( .A(n3895), .B(n23450), .Y(n23451) );
  INVX1 U5307 ( .A(n19887), .Y(n20059) );
  INVX1 U5308 ( .A(n20156), .Y(n20083) );
  INVXL U5309 ( .A(n5465), .Y(n23556) );
  NAND3X2 U5310 ( .A(n4198), .B(n5436), .C(n18973), .Y(n23561) );
  INVX1 U5311 ( .A(n3084), .Y(n3859) );
  AOI21X1 U5312 ( .A0(n20018), .A1(n19763), .B0(n19762), .Y(n19887) );
  NAND2X1 U5313 ( .A(n3357), .B(n17424), .Y(n17426) );
  INVX1 U5314 ( .A(n20808), .Y(n20752) );
  XNOR2X1 U5315 ( .A(n10967), .B(n10966), .Y(n23541) );
  NAND2XL U5316 ( .A(n3357), .B(n17451), .Y(n17454) );
  NOR2BX2 U5317 ( .AN(n23529), .B(n3033), .Y(n23512) );
  AOI21X1 U5318 ( .A0(n8403), .A1(n8643), .B0(n8642), .Y(n8644) );
  NAND2XL U5319 ( .A(n3357), .B(n20735), .Y(n6045) );
  AOI21XL U5320 ( .A0(n15261), .A1(n15657), .B0(n15370), .Y(n15371) );
  NAND2X1 U5321 ( .A(n3357), .B(n17444), .Y(n17447) );
  NAND3X1 U5322 ( .A(n23456), .B(n6033), .C(n23515), .Y(n18975) );
  NAND2X1 U5323 ( .A(n5100), .B(n20856), .Y(n10743) );
  NAND2X1 U5324 ( .A(n5100), .B(n10740), .Y(n10742) );
  NOR2X2 U5325 ( .A(n3446), .B(n3344), .Y(n4652) );
  NAND2X1 U5326 ( .A(n5100), .B(n20892), .Y(n3456) );
  INVX1 U5327 ( .A(n4001), .Y(n17456) );
  AOI21X1 U5328 ( .A0(n19907), .A1(n19983), .B0(n19906), .Y(n19908) );
  OR2XL U5329 ( .A(n19702), .B(n19701), .Y(n20069) );
  NAND3XL U5330 ( .A(n18973), .B(n6024), .C(n24250), .Y(n18974) );
  AOI21X1 U5331 ( .A0(n15527), .A1(n15604), .B0(n15526), .Y(n15528) );
  NOR3X2 U5332 ( .A(n17359), .B(n5699), .C(n3931), .Y(n3339) );
  NAND2X1 U5333 ( .A(n3304), .B(n10637), .Y(n10642) );
  NOR2X1 U5334 ( .A(n3931), .B(n5699), .Y(n3864) );
  INVX1 U5335 ( .A(n6024), .Y(n4395) );
  INVX1 U5336 ( .A(n21043), .Y(n20669) );
  XOR2X1 U5337 ( .A(n19062), .B(n20954), .Y(n20956) );
  NAND2X1 U5338 ( .A(n5719), .B(n23641), .Y(n5698) );
  NAND2X1 U5339 ( .A(n21836), .B(n22105), .Y(n21838) );
  INVX1 U5340 ( .A(n23589), .Y(n23590) );
  NAND2X1 U5341 ( .A(n20982), .B(n20980), .Y(n5273) );
  NOR2X1 U5342 ( .A(n8831), .B(n8835), .Y(n8826) );
  NAND3BX2 U5343 ( .AN(n3989), .B(n3987), .C(n3986), .Y(n20671) );
  NAND2X1 U5344 ( .A(n15447), .B(n15446), .Y(n15494) );
  NAND2XL U5345 ( .A(n8649), .B(n8648), .Y(n8764) );
  INVX1 U5346 ( .A(n20348), .Y(n20360) );
  NAND2XL U5347 ( .A(n8647), .B(n8646), .Y(n8920) );
  INVXL U5348 ( .A(n22198), .Y(n22193) );
  NAND2X1 U5349 ( .A(n15525), .B(n15524), .Y(n15615) );
  NAND2X1 U5350 ( .A(n15563), .B(n15562), .Y(n15593) );
  XOR2X2 U5351 ( .A(n4021), .B(n12889), .Y(n21019) );
  NAND2X1 U5352 ( .A(n15394), .B(n15393), .Y(n15670) );
  NAND2X2 U5353 ( .A(n18422), .B(n18918), .Y(n3431) );
  INVX1 U5354 ( .A(n10998), .Y(n11353) );
  NAND2X1 U5355 ( .A(n15565), .B(n15564), .Y(n15626) );
  NAND2X1 U5356 ( .A(n19777), .B(n19776), .Y(n19893) );
  NAND2X1 U5357 ( .A(n15396), .B(n15395), .Y(n15513) );
  NAND2X1 U5358 ( .A(n8776), .B(n8775), .Y(n8865) );
  NAND2X1 U5359 ( .A(n19775), .B(n19774), .Y(n20049) );
  NAND2XL U5360 ( .A(n15443), .B(n15442), .Y(n15504) );
  NAND2XL U5361 ( .A(n8694), .B(n8693), .Y(n8755) );
  OAI2BB1X1 U5362 ( .A0N(n5681), .A1N(n3781), .B0(n5683), .Y(n5682) );
  NOR2X2 U5363 ( .A(n12921), .B(n12929), .Y(n3347) );
  INVX1 U5364 ( .A(n23481), .Y(n4160) );
  NAND2XL U5365 ( .A(n19823), .B(n19822), .Y(n19884) );
  CLKINVX3 U5366 ( .A(n17425), .Y(n17421) );
  NAND2X1 U5367 ( .A(n19942), .B(n19941), .Y(n19972) );
  AOI21XL U5368 ( .A0(n14674), .A1(n14535), .B0(n14534), .Y(n14536) );
  BUFX16 U5369 ( .A(n3469), .Y(n3415) );
  AOI21XL U5370 ( .A0(n14674), .A1(n14543), .B0(n14542), .Y(n14544) );
  INVX1 U5371 ( .A(n22114), .Y(n22099) );
  OR2X1 U5372 ( .A(n15359), .B(n15187), .Y(n15189) );
  AOI21X1 U5373 ( .A0(n15556), .A1(n23955), .B0(n15573), .Y(n15555) );
  INVX1 U5374 ( .A(n20816), .Y(n20817) );
  OR2X1 U5375 ( .A(n8506), .B(n8614), .Y(n8508) );
  NOR2X1 U5376 ( .A(n10729), .B(n20896), .Y(n7452) );
  NAND2X1 U5377 ( .A(n19944), .B(n19943), .Y(n20005) );
  INVX1 U5378 ( .A(n20278), .Y(n20858) );
  NOR2X2 U5379 ( .A(n20893), .B(n20896), .Y(n3536) );
  INVXL U5380 ( .A(n20618), .Y(n20619) );
  NAND2X1 U5381 ( .A(n8295), .B(n8769), .Y(n8771) );
  OR2X2 U5382 ( .A(n21826), .B(n21825), .Y(n6202) );
  NAND2X1 U5383 ( .A(n15046), .B(n15539), .Y(n15541) );
  OR2X1 U5384 ( .A(n19748), .B(n19717), .Y(n19719) );
  INVX1 U5385 ( .A(n12973), .Y(n12975) );
  NAND2BX1 U5386 ( .AN(n12810), .B(n12865), .Y(n4051) );
  NAND2X1 U5387 ( .A(n8295), .B(n8785), .Y(n8787) );
  NAND2X1 U5388 ( .A(n10505), .B(n4611), .Y(n10603) );
  AOI21X1 U5389 ( .A0(n10608), .A1(n4611), .B0(n10470), .Y(n10604) );
  OR2X1 U5390 ( .A(n21814), .B(n21813), .Y(n21792) );
  NAND2XL U5391 ( .A(n19424), .B(n19919), .Y(n19921) );
  NAND2X1 U5392 ( .A(n22002), .B(n22001), .Y(n22031) );
  NOR2X1 U5393 ( .A(n19553), .B(n19807), .Y(n19838) );
  INVXL U5394 ( .A(n22027), .Y(n22066) );
  NOR2X1 U5395 ( .A(n15244), .B(n3090), .Y(n15518) );
  NOR2X1 U5396 ( .A(n8476), .B(n3154), .Y(n8709) );
  AND2X2 U5397 ( .A(n10224), .B(n10223), .Y(n4605) );
  INVXL U5398 ( .A(n10612), .Y(n10504) );
  NAND2X1 U5399 ( .A(n14526), .B(n14525), .Y(n14527) );
  AOI2BB2X1 U5400 ( .B0(n8322), .B1(n3157), .A0N(n3157), .A1N(n8463), .Y(n8476) );
  NAND2X1 U5401 ( .A(n14556), .B(n14555), .Y(n14557) );
  OR2XL U5402 ( .A(n21753), .B(n21787), .Y(n21755) );
  NAND2X1 U5403 ( .A(n22006), .B(n22005), .Y(n22072) );
  NOR2X1 U5404 ( .A(n11363), .B(n11370), .Y(n11386) );
  NAND2BX1 U5405 ( .AN(n10477), .B(n5219), .Y(n4364) );
  NAND2XL U5406 ( .A(n5621), .B(n7256), .Y(n7007) );
  INVX1 U5407 ( .A(n13981), .Y(n13647) );
  NAND2BX1 U5408 ( .AN(n15318), .B(n15289), .Y(n15350) );
  NAND2X1 U5409 ( .A(n12978), .B(n12853), .Y(n12855) );
  AOI2BB2X1 U5410 ( .B0(n19451), .B1(n19542), .A0N(n19542), .A1N(n19741), .Y(
        n19553) );
  INVX1 U5411 ( .A(n10195), .Y(n10227) );
  AOI21X1 U5412 ( .A0(n14397), .A1(n3152), .B0(n4483), .Y(n4482) );
  CLKINVX3 U5413 ( .A(n3154), .Y(n3086) );
  AOI2BB2X1 U5414 ( .B0(n19714), .B1(n19542), .A0N(n19542), .A1N(n19713), .Y(
        n19782) );
  NAND2X1 U5415 ( .A(n17233), .B(n17232), .Y(n17234) );
  INVX1 U5416 ( .A(n17216), .Y(n17250) );
  OR2XL U5417 ( .A(n21787), .B(n21786), .Y(n21789) );
  OR2XL U5418 ( .A(n21787), .B(n21772), .Y(n21774) );
  AOI2BB2XL U5419 ( .B0(n3036), .B1(n19712), .A0N(n3036), .A1N(n19711), .Y(
        n19783) );
  NAND2XL U5420 ( .A(n3156), .B(n3167), .Y(n15318) );
  INVX1 U5421 ( .A(n10607), .Y(n10615) );
  OAI21XL U5422 ( .A0(n3163), .A1(n3324), .B0(n3323), .Y(n10443) );
  INVX1 U5423 ( .A(n17207), .Y(n17209) );
  NAND2X1 U5424 ( .A(n21506), .B(n21979), .Y(n21981) );
  ADDFHX2 U5425 ( .A(n9412), .B(n9411), .CI(n9410), .CO(n10130), .S(n10129) );
  INVX1 U5426 ( .A(n17239), .Y(n3158) );
  AOI21XL U5427 ( .A0(n17312), .A1(n17328), .B0(n17327), .Y(n17329) );
  NAND2X1 U5428 ( .A(n3035), .B(n3039), .Y(n19467) );
  NAND2XL U5429 ( .A(n10437), .B(n3322), .Y(n3323) );
  INVXL U5430 ( .A(n12895), .Y(n3886) );
  INVX1 U5431 ( .A(n10469), .Y(n3305) );
  INVXL U5432 ( .A(n18834), .Y(n18836) );
  NOR2X2 U5433 ( .A(n18393), .B(n18392), .Y(n18727) );
  INVXL U5434 ( .A(n9764), .Y(n3277) );
  NAND2X1 U5435 ( .A(n21506), .B(n21974), .Y(n21976) );
  INVXL U5436 ( .A(n20646), .Y(n20636) );
  NOR2X1 U5437 ( .A(n21846), .B(n3171), .Y(n21979) );
  NAND2X1 U5438 ( .A(n3162), .B(n3092), .Y(n8337) );
  INVX1 U5439 ( .A(n18322), .Y(n4179) );
  AOI21X1 U5440 ( .A0(n4236), .A1(n4235), .B0(n4233), .Y(n4232) );
  AND2X1 U5441 ( .A(n21855), .B(n21793), .Y(n21984) );
  NAND2XL U5442 ( .A(n3037), .B(n21707), .Y(n21720) );
  NAND2X1 U5443 ( .A(n18690), .B(n3000), .Y(n18692) );
  INVX1 U5444 ( .A(n17315), .Y(n4943) );
  AOI21XL U5445 ( .A0(n12808), .A1(n12794), .B0(n12793), .Y(n12825) );
  NOR2X1 U5446 ( .A(n21839), .B(n3171), .Y(n21974) );
  INVX4 U5447 ( .A(n4591), .Y(n3162) );
  ADDFHX1 U5448 ( .A(n18385), .B(n18384), .CI(n18383), .CO(n18392), .S(n18322)
         );
  INVXL U5449 ( .A(n7020), .Y(n7022) );
  INVXL U5450 ( .A(n12856), .Y(n12837) );
  NAND2X1 U5451 ( .A(n4231), .B(n4230), .Y(n4229) );
  NAND2X2 U5452 ( .A(n12497), .B(n12496), .Y(n12895) );
  ADDFHX1 U5453 ( .A(n13744), .B(n13743), .CI(n13742), .CO(n13802), .S(n13820)
         );
  NAND2XL U5454 ( .A(n3163), .B(n3324), .Y(n3322) );
  INVX1 U5455 ( .A(n3280), .Y(n3278) );
  NAND2XL U5456 ( .A(n9691), .B(n9692), .Y(n6067) );
  AOI22XL U5457 ( .A0(n21742), .A1(n3171), .B0(n21741), .B1(n3037), .Y(n21877)
         );
  NOR2X1 U5458 ( .A(n21742), .B(n3171), .Y(n22011) );
  NAND2XL U5459 ( .A(n9414), .B(n9415), .Y(n5307) );
  INVX1 U5460 ( .A(n7443), .Y(n3168) );
  OAI21X1 U5461 ( .A0(n7792), .A1(n7791), .B0(n7790), .Y(n7819) );
  INVX1 U5462 ( .A(n21696), .Y(n21783) );
  NAND2X1 U5463 ( .A(n3473), .B(n3474), .Y(n3472) );
  NAND2X1 U5464 ( .A(n3093), .B(n3097), .Y(n18318) );
  CLKINVX3 U5465 ( .A(n3171), .Y(n3037) );
  AOI2BB2X1 U5466 ( .B0(n21769), .B1(n3096), .A0N(n3096), .A1N(n21768), .Y(
        n21839) );
  XNOR2X1 U5467 ( .A(n8232), .B(n8231), .Y(n4591) );
  NOR2X2 U5468 ( .A(n12936), .B(n12933), .Y(n12873) );
  ADDFHX2 U5469 ( .A(n12474), .B(n12473), .CI(n12472), .CO(n12496), .S(n12495)
         );
  INVX1 U5470 ( .A(n10438), .Y(n3324) );
  ADDFHX1 U5471 ( .A(n10436), .B(n10435), .CI(n10434), .CO(n10441), .S(n10444)
         );
  INVX1 U5472 ( .A(n18941), .Y(n18947) );
  ADDFHX2 U5473 ( .A(n11866), .B(n11865), .CI(n11864), .CO(n12498), .S(n12497)
         );
  NAND2XL U5474 ( .A(n7005), .B(n7255), .Y(n7006) );
  NAND2X1 U5475 ( .A(n10502), .B(n10501), .Y(n10551) );
  INVX1 U5476 ( .A(n18848), .Y(n18851) );
  OAI21XL U5477 ( .A0(n12688), .A1(n12689), .B0(n12687), .Y(n4932) );
  NOR2X2 U5478 ( .A(n17348), .B(n17326), .Y(n17122) );
  NOR2X1 U5479 ( .A(M6_mult_x_15_n483), .B(M6_mult_x_15_n490), .Y(n11357) );
  AOI21X2 U5480 ( .A0(n7728), .A1(n7727), .B0(n7726), .Y(n7792) );
  NOR2X1 U5481 ( .A(n7788), .B(n7791), .Y(n7814) );
  INVX4 U5482 ( .A(n4618), .Y(n3171) );
  INVX1 U5483 ( .A(n18316), .Y(n3093) );
  INVX1 U5484 ( .A(n17115), .Y(n5057) );
  INVX1 U5485 ( .A(n15015), .Y(n4458) );
  NOR2X1 U5486 ( .A(n10978), .B(n10973), .Y(n11005) );
  NAND2X1 U5487 ( .A(n24431), .B(n15027), .Y(n15033) );
  INVX1 U5488 ( .A(n18678), .Y(n4251) );
  INVXL U5489 ( .A(n12416), .Y(n4981) );
  ADDFHX2 U5490 ( .A(n16298), .B(n16297), .CI(n16296), .CO(n16865), .S(n16863)
         );
  ADDFHX1 U5491 ( .A(n10304), .B(n10303), .CI(n10302), .CO(n10438), .S(n10317)
         );
  INVXL U5492 ( .A(n9522), .Y(n5521) );
  INVX1 U5493 ( .A(n17116), .Y(n5686) );
  INVX4 U5494 ( .A(n15004), .Y(n15289) );
  ADDFHX1 U5495 ( .A(n10086), .B(n10085), .CI(n10084), .CO(n10065), .S(n10101)
         );
  ADDFHX2 U5496 ( .A(n12094), .B(n12093), .CI(n12092), .CO(n12087), .S(n12112)
         );
  NAND2BX1 U5497 ( .AN(n12722), .B(n12871), .Y(n12788) );
  ADDFHX2 U5498 ( .A(n16138), .B(n16137), .CI(n16136), .CO(n16189), .S(n16152)
         );
  NAND2X1 U5499 ( .A(n8280), .B(n8285), .Y(n8282) );
  INVX1 U5500 ( .A(n17113), .Y(n5056) );
  ADDFHX1 U5501 ( .A(n17988), .B(n17987), .CI(n17986), .CO(n18319), .S(n18316)
         );
  ADDFHX2 U5502 ( .A(n11904), .B(n11903), .CI(n11902), .CO(n12508), .S(n12506)
         );
  AND2X2 U5503 ( .A(n7764), .B(n7762), .Y(n4609) );
  INVX1 U5504 ( .A(n18959), .Y(n18961) );
  AOI21X2 U5505 ( .A0(n17592), .A1(n5022), .B0(n3427), .Y(n5865) );
  OAI21X1 U5506 ( .A0(n11824), .A1(n11825), .B0(n11823), .Y(n4024) );
  NOR2X1 U5507 ( .A(M6_mult_x_15_n463), .B(M6_mult_x_15_n468), .Y(n10978) );
  NAND2BXL U5508 ( .AN(n16774), .B(n5544), .Y(n16505) );
  NOR2X1 U5509 ( .A(n18695), .B(n18696), .Y(n18942) );
  INVXL U5510 ( .A(n16773), .Y(n5544) );
  INVXL U5511 ( .A(n16953), .Y(n5830) );
  CLKINVX2 U5512 ( .A(n6731), .Y(n5636) );
  INVX1 U5513 ( .A(n6730), .Y(n3572) );
  INVXL U5514 ( .A(n16765), .Y(n3945) );
  INVXL U5515 ( .A(n12481), .Y(n3907) );
  NOR2X1 U5516 ( .A(n23870), .B(n8222), .Y(n8228) );
  NOR2X1 U5517 ( .A(n23760), .B(n8233), .Y(n8231) );
  OAI21XL U5518 ( .A0(n17843), .A1(n17844), .B0(n17842), .Y(n5901) );
  XOR3X2 U5519 ( .A(n17644), .B(n17643), .C(n17642), .Y(n17647) );
  XOR2X2 U5520 ( .A(n3706), .B(n16432), .Y(n16450) );
  NAND2X1 U5521 ( .A(n6078), .B(n6077), .Y(n17570) );
  XOR2X1 U5522 ( .A(n4961), .B(n12386), .Y(n3997) );
  OAI21XL U5523 ( .A0(n17003), .A1(n17004), .B0(n3954), .Y(n4100) );
  NAND2XL U5524 ( .A(n12476), .B(n5775), .Y(n5773) );
  NOR2X1 U5525 ( .A(n23179), .B(n23178), .Y(n8213) );
  OAI2BB1X1 U5526 ( .A0N(n17067), .A1N(n17065), .B0(n5094), .Y(n17130) );
  INVX1 U5527 ( .A(n23180), .Y(n8275) );
  OAI2BB1X1 U5528 ( .A0N(n11785), .A1N(n4863), .B0(n4862), .Y(n11870) );
  OAI22XL U5529 ( .A0(n15538), .A1(n3101), .B0(n15008), .B1(n15537), .Y(n15560) );
  INVX1 U5530 ( .A(n16434), .Y(n3705) );
  OAI21X1 U5531 ( .A0(n16018), .A1(n16019), .B0(n16017), .Y(n3341) );
  INVXL U5532 ( .A(n4881), .Y(n4004) );
  ADDFHX2 U5533 ( .A(n16097), .B(n16096), .CI(n16095), .CO(n16081), .S(n16804)
         );
  XOR2X1 U5534 ( .A(n11720), .B(n11719), .Y(n4430) );
  ADDFHX2 U5535 ( .A(n16295), .B(n16294), .CI(n16293), .CO(n16862), .S(n16860)
         );
  OAI2BB1X1 U5536 ( .A0N(n12444), .A1N(n12443), .B0(n5404), .Y(n12481) );
  ADDFHX1 U5537 ( .A(n12459), .B(n12458), .CI(n12457), .CO(n12477), .S(n12468)
         );
  NAND2X1 U5538 ( .A(n21488), .B(n21487), .Y(n21489) );
  ADDFHX2 U5539 ( .A(n17984), .B(n17983), .CI(n17982), .CO(n17957), .S(n17986)
         );
  NOR2BXL U5540 ( .AN(n24043), .B(n24042), .Y(n24045) );
  ADDFHX2 U5541 ( .A(n6812), .B(n6810), .CI(n6811), .CO(n6907), .S(n6906) );
  INVXL U5542 ( .A(n17686), .Y(n4314) );
  ADDFHX1 U5543 ( .A(n6389), .B(n6388), .CI(n6387), .CO(n6731), .S(n6730) );
  INVXL U5544 ( .A(n3269), .Y(n3266) );
  NAND2XL U5545 ( .A(n3287), .B(n3288), .Y(n3299) );
  OAI21X1 U5546 ( .A0(n21450), .A1(n21453), .B0(n21451), .Y(n21483) );
  OAI2BB1X1 U5547 ( .A0N(n5414), .A1N(n4075), .B0(n5412), .Y(n12626) );
  NAND2XL U5548 ( .A(n12175), .B(n4486), .Y(n4020) );
  XOR2X1 U5549 ( .A(n12134), .B(n3388), .Y(n3387) );
  INVX1 U5550 ( .A(n21501), .Y(n21503) );
  INVXL U5551 ( .A(n3388), .Y(n3385) );
  INVX1 U5552 ( .A(n23210), .Y(n19363) );
  OAI22X1 U5553 ( .A0(n8773), .A1(n3017), .B0(n3040), .B1(n8772), .Y(n8775) );
  XOR3X4 U5554 ( .A(n18337), .B(n18336), .C(n18335), .Y(n18358) );
  OAI22XL U5555 ( .A0(n15553), .A1(n3101), .B0(n15558), .B1(n15552), .Y(n15566) );
  OAI22X1 U5556 ( .A0(n8789), .A1(n3017), .B0(n3040), .B1(n8788), .Y(n8810) );
  OAI21X1 U5557 ( .A0(n15558), .A1(n14945), .B0(n14944), .Y(n23163) );
  NAND2BX1 U5558 ( .AN(n18264), .B(n3358), .Y(n18267) );
  XNOR2X1 U5559 ( .A(n3352), .B(n4864), .Y(n4863) );
  OAI22X1 U5560 ( .A0(n10541), .A1(n25885), .B0(n10540), .B1(n3174), .Y(n10549) );
  NAND2X1 U5561 ( .A(n10541), .B(n3174), .Y(n5751) );
  INVX1 U5562 ( .A(n9504), .Y(n3099) );
  NAND2X1 U5563 ( .A(n15190), .B(n14950), .Y(n14916) );
  NAND2X1 U5564 ( .A(n15190), .B(n14954), .Y(n14914) );
  NAND2X1 U5565 ( .A(n15190), .B(n14951), .Y(n14952) );
  OAI22X1 U5566 ( .A0(n19923), .A1(n3100), .B0(n3041), .B1(n19922), .Y(n19941)
         );
  INVX1 U5567 ( .A(n12431), .Y(n3651) );
  OAI22X1 U5568 ( .A0(n19918), .A1(n3100), .B0(n3041), .B1(n19917), .Y(n19939)
         );
  ADDFHX1 U5569 ( .A(n11822), .B(n11821), .CI(n11820), .CO(n11860), .S(n12475)
         );
  NOR2X1 U5570 ( .A(n3271), .B(n3270), .Y(n3269) );
  OAI2BB1XL U5571 ( .A0N(n5517), .A1N(n6062), .B0(n6060), .Y(n9300) );
  CLKINVX2 U5572 ( .A(n12113), .Y(n3474) );
  OAI22X1 U5573 ( .A0(n19933), .A1(n3100), .B0(n3041), .B1(n19932), .Y(n19945)
         );
  NAND2X1 U5574 ( .A(n8482), .B(n8196), .Y(n8197) );
  NAND2X1 U5575 ( .A(n8482), .B(n8185), .Y(n8186) );
  NAND2BXL U5576 ( .AN(n16053), .B(n3633), .Y(n3632) );
  ADDFHX2 U5577 ( .A(n16817), .B(n16816), .CI(n16815), .CO(n16810), .S(n16834)
         );
  NAND2BXL U5578 ( .AN(n13792), .B(n13258), .Y(n5487) );
  ADDFHX1 U5579 ( .A(n16996), .B(n16995), .CI(n16994), .CO(n17003), .S(n17021)
         );
  NAND2XL U5580 ( .A(n4194), .B(n18362), .Y(n4091) );
  NAND2XL U5581 ( .A(n23413), .B(n21493), .Y(n21497) );
  NOR2X1 U5582 ( .A(n23230), .B(n21485), .Y(n21501) );
  NAND2X1 U5583 ( .A(n23230), .B(n21485), .Y(n21502) );
  OAI2BB1XL U5584 ( .A0N(n4045), .A1N(n12581), .B0(n4044), .Y(n12690) );
  ADDFHX1 U5585 ( .A(n17684), .B(n17683), .CI(n17682), .CO(n17726), .S(n18335)
         );
  NOR2X1 U5586 ( .A(n23420), .B(n21444), .Y(n21450) );
  ADDFHX1 U5587 ( .A(n18349), .B(n18348), .CI(n18347), .CO(n18375), .S(n18368)
         );
  NOR2X1 U5588 ( .A(n6084), .B(n6083), .Y(n6082) );
  INVX1 U5589 ( .A(n23121), .Y(n21485) );
  ADDFHX2 U5590 ( .A(n11682), .B(n11681), .CI(n11680), .CO(n11692), .S(n11790)
         );
  OR2XL U5591 ( .A(n7179), .B(n7178), .Y(n3544) );
  NOR2XL U5592 ( .A(n10668), .B(n10667), .Y(n10669) );
  OAI21XL U5593 ( .A0(n7141), .A1(n7140), .B0(n7139), .Y(n5564) );
  ADDFHX1 U5594 ( .A(n12146), .B(n12145), .CI(n12144), .CO(n12158), .S(n12176)
         );
  XOR2X1 U5595 ( .A(n6498), .B(n5633), .Y(n6519) );
  NAND2BXL U5596 ( .AN(n5805), .B(n16428), .Y(n5803) );
  OAI21X1 U5597 ( .A0(n21519), .A1(n21428), .B0(n21427), .Y(n23124) );
  OAI2BB1X1 U5598 ( .A0N(n17591), .A1N(n5923), .B0(n5922), .Y(n17598) );
  ADDFHX1 U5599 ( .A(n6336), .B(n6335), .CI(n6334), .CO(n6806), .S(n6385) );
  NAND2BXL U5600 ( .AN(n3846), .B(n5980), .Y(n5979) );
  AND2X1 U5601 ( .A(n19042), .B(n19041), .Y(n22481) );
  INVXL U5602 ( .A(n3929), .Y(n3928) );
  OR2X2 U5603 ( .A(n18724), .B(n18723), .Y(n18726) );
  ADDFHX1 U5604 ( .A(n16134), .B(n16133), .CI(n16132), .CO(n16159), .S(n16148)
         );
  OAI21X1 U5605 ( .A0(n17536), .A1(n18168), .B0(n3412), .Y(n17663) );
  INVXL U5606 ( .A(n16114), .Y(n3685) );
  OAI22XL U5607 ( .A0(n12759), .A1(n12700), .B0(n12760), .B1(n12713), .Y(
        n12709) );
  OAI21XL U5608 ( .A0(n3106), .A1(n3107), .B0(n3967), .Y(n12708) );
  OAI22X1 U5609 ( .A0(n12759), .A1(n11984), .B0(n12760), .B1(n12637), .Y(
        n12613) );
  OAI22X1 U5610 ( .A0(n12635), .A1(n11792), .B0(n12513), .B1(n4512), .Y(n11833) );
  INVX8 U5611 ( .A(n8161), .Y(n3017) );
  INVX1 U5612 ( .A(n3564), .Y(n3561) );
  OAI22X1 U5613 ( .A0(n16701), .A1(n16051), .B0(n16699), .B1(n16050), .Y(
        n16090) );
  XOR2XL U5614 ( .A(n17624), .B(n6125), .Y(n17633) );
  NAND3XL U5615 ( .A(n9153), .B(n9152), .C(n14452), .Y(n10693) );
  XOR2X1 U5616 ( .A(n17181), .B(n17403), .Y(n17196) );
  OAI22X1 U5617 ( .A0(n18083), .A1(n17942), .B0(n18429), .B1(n17879), .Y(n4394) );
  OAI22X1 U5618 ( .A0(n3102), .A1(n3780), .B0(n16332), .B1(n16088), .Y(n16105)
         );
  OAI21X1 U5619 ( .A0(n16518), .A1(n16475), .B0(n3789), .Y(n16529) );
  OAI22X1 U5620 ( .A0(n3102), .A1(n16009), .B0(n16332), .B1(n15964), .Y(n16053) );
  OAI21X2 U5621 ( .A0(n22506), .A1(n11081), .B0(n11080), .Y(n11082) );
  OAI22X1 U5622 ( .A0(n18659), .A1(n17742), .B0(n17832), .B1(n17777), .Y(
        n17788) );
  INVX1 U5623 ( .A(n17074), .Y(n5066) );
  NAND2X1 U5624 ( .A(n3414), .B(n3413), .Y(n3412) );
  XNOR2X1 U5625 ( .A(n7830), .B(n25872), .Y(n7831) );
  NAND2BXL U5626 ( .AN(n17655), .B(n5896), .Y(n5768) );
  OR2X1 U5627 ( .A(n17045), .B(n17099), .Y(n5825) );
  NAND2XL U5628 ( .A(n5893), .B(n18541), .Y(n5894) );
  XOR2X1 U5629 ( .A(n11588), .B(n13010), .Y(n11616) );
  INVXL U5630 ( .A(n5415), .Y(n3841) );
  OAI21X1 U5631 ( .A0(n16381), .A1(n16704), .B0(n3702), .Y(n16439) );
  AOI21X1 U5632 ( .A0(n21085), .A1(n11069), .B0(n11068), .Y(n22506) );
  NAND2XL U5633 ( .A(n2992), .B(n3044), .Y(n3698) );
  OR2XL U5634 ( .A(n6013), .B(n16965), .Y(n6012) );
  INVX4 U5635 ( .A(n21429), .Y(n3020) );
  OAI22X1 U5636 ( .A0(n16686), .A1(n16685), .B0(n16684), .B1(n16475), .Y(
        n16694) );
  INVX1 U5637 ( .A(n18242), .Y(n3414) );
  OAI22XL U5638 ( .A0(n6501), .A1(n6845), .B0(n6497), .B1(n6843), .Y(n6520) );
  INVXL U5639 ( .A(n13769), .Y(n13100) );
  OAI211X1 U5640 ( .A0(n24001), .A1(n25243), .B0(n9095), .C0(n11514), .Y(
        M2_b_0_) );
  XNOR2X1 U5641 ( .A(n25884), .B(n5430), .Y(n11743) );
  OAI2BB1X1 U5642 ( .A0N(n17832), .A1N(n18666), .B0(n25883), .Y(n18671) );
  XOR2X1 U5643 ( .A(n5677), .B(n3048), .Y(n5061) );
  XNOR2X1 U5644 ( .A(n5677), .B(n3201), .Y(n16868) );
  CLKINVX3 U5645 ( .A(n7040), .Y(n6366) );
  AND2X2 U5646 ( .A(n17148), .B(n17147), .Y(n17149) );
  XOR2X2 U5647 ( .A(n4888), .B(n3210), .Y(n17501) );
  OR2XL U5648 ( .A(n11648), .B(n12222), .Y(n5324) );
  BUFX3 U5649 ( .A(M1_a_4_), .Y(n25865) );
  NAND2XL U5650 ( .A(n4566), .B(learning_rate[2]), .Y(n4551) );
  NAND2BX1 U5651 ( .AN(n14700), .B(n14698), .Y(n14449) );
  OAI21XL U5652 ( .A0(n19193), .A1(n19192), .B0(n19191), .Y(n19194) );
  NOR2BX1 U5653 ( .AN(n3110), .B(n12995), .Y(n11751) );
  OAI21XL U5654 ( .A0(n19148), .A1(n19147), .B0(n19146), .Y(n19196) );
  XNOR2X1 U5655 ( .A(n12732), .B(n12560), .Y(n11985) );
  CLKBUFX2 U5656 ( .A(M1_a_8_), .Y(n4565) );
  XOR2X1 U5657 ( .A(n12701), .B(n3191), .Y(n3883) );
  NAND2XL U5658 ( .A(n15946), .B(n15947), .Y(n16570) );
  BUFX12 U5659 ( .A(M3_mult_x_15_b_11_), .Y(n3190) );
  AOI21X1 U5660 ( .A0(n19190), .A1(n19189), .B0(n19188), .Y(n19191) );
  AOI21X1 U5661 ( .A0(n19280), .A1(n19239), .B0(n19279), .Y(n19281) );
  AOI22XL U5662 ( .A0(n22486), .A1(sigma12[21]), .B0(n25750), .B1(sigma11[21]), 
        .Y(n25751) );
  BUFX12 U5663 ( .A(M3_mult_x_15_b_17_), .Y(n3201) );
  INVX8 U5664 ( .A(n16873), .Y(n3203) );
  NOR2X1 U5665 ( .A(n8666), .B(n8263), .Y(n8008) );
  NOR2X1 U5666 ( .A(n8681), .B(n8236), .Y(n8014) );
  AND2X2 U5667 ( .A(n3111), .B(data[126]), .Y(n17155) );
  INVX4 U5668 ( .A(n5729), .Y(n15968) );
  BUFX3 U5669 ( .A(n17459), .Y(n25750) );
  AND2X2 U5670 ( .A(n3111), .B(data[94]), .Y(n18737) );
  INVXL U5671 ( .A(M3_mult_x_15_b_1_), .Y(n11697) );
  NOR2XL U5672 ( .A(n8169), .B(n8207), .Y(n8097) );
  OR2XL U5673 ( .A(n9109), .B(n3218), .Y(n11070) );
  OR2XL U5674 ( .A(n11071), .B(n3218), .Y(n11072) );
  NOR2XL U5675 ( .A(n4527), .B(n4526), .Y(n4525) );
  NAND2X1 U5676 ( .A(n21272), .B(n21246), .Y(n21259) );
  NOR2X1 U5677 ( .A(n19532), .B(n19486), .Y(n19142) );
  NOR2X1 U5678 ( .A(n19802), .B(n19364), .Y(n19165) );
  INVX1 U5679 ( .A(n7569), .Y(n7550) );
  INVX1 U5680 ( .A(n8254), .Y(n8326) );
  NOR2X1 U5681 ( .A(n14734), .B(n14795), .Y(n14740) );
  AOI21XL U5682 ( .A0(n21285), .A1(n21284), .B0(n21283), .Y(n21286) );
  NOR2X1 U5683 ( .A(n19841), .B(n19435), .Y(n19201) );
  NAND2X2 U5684 ( .A(n4518), .B(n6090), .Y(M4_a_7_) );
  OAI2BB1X1 U5685 ( .A0N(learning_rate[9]), .A1N(in_valid_t), .B0(n6163), .Y(
        n3333) );
  BUFX4 U5686 ( .A(n11488), .Y(M3_mult_x_15_b_6_) );
  INVX1 U5687 ( .A(n25206), .Y(n20353) );
  INVX1 U5688 ( .A(n8408), .Y(n8420) );
  INVX4 U5689 ( .A(n20373), .Y(n25743) );
  INVX1 U5690 ( .A(n5158), .Y(n4250) );
  CLKINVX3 U5691 ( .A(M0_a_2_), .Y(n3591) );
  BUFX2 U5692 ( .A(n25785), .Y(n25763) );
  OAI2BB1X1 U5693 ( .A0N(y10[25]), .A1N(n3224), .B0(n7398), .Y(n7856) );
  INVX4 U5694 ( .A(n3584), .Y(n25874) );
  AOI22X1 U5695 ( .A0(n5770), .A1(data[71]), .B0(in_valid_t), .B1(w2[39]), .Y(
        n4518) );
  NOR2X1 U5696 ( .A(n19255), .B(n19325), .Y(n19258) );
  NOR2X1 U5697 ( .A(n19932), .B(n19427), .Y(n19254) );
  NAND4X1 U5698 ( .A(n7935), .B(n7934), .C(n7933), .D(n7932), .Y(n8355) );
  AND2XL U5699 ( .A(n5015), .B(data[90]), .Y(n18748) );
  INVX4 U5700 ( .A(n3117), .Y(n3051) );
  OAI21X1 U5701 ( .A0(n7382), .A1(n26000), .B0(n6234), .Y(M0_a_2_) );
  NAND2XL U5702 ( .A(n5480), .B(sigma11[2]), .Y(n5049) );
  INVX1 U5703 ( .A(n19485), .Y(n19508) );
  NAND2XL U5704 ( .A(n5480), .B(sigma11[8]), .Y(n6089) );
  INVX4 U5705 ( .A(n3117), .Y(n3023) );
  CLKINVX8 U5706 ( .A(n3117), .Y(n3052) );
  NOR2X1 U5707 ( .A(n21337), .B(n21514), .Y(n21301) );
  NOR2X1 U5708 ( .A(n21350), .B(n21509), .Y(n21313) );
  NAND2X1 U5709 ( .A(n8104), .B(y20[25]), .Y(n8081) );
  BUFX3 U5710 ( .A(n11147), .Y(n11062) );
  CLKINVX3 U5711 ( .A(n22490), .Y(n3053) );
  INVX1 U5712 ( .A(n15175), .Y(n15206) );
  NAND2X1 U5713 ( .A(n3120), .B(y20[24]), .Y(n8077) );
  AOI21XL U5714 ( .A0(n21166), .A1(sigma12[9]), .B0(n5730), .Y(n4101) );
  NAND2XL U5715 ( .A(n21166), .B(target_temp[30]), .Y(n11550) );
  XOR2X1 U5716 ( .A(n3058), .B(n21059), .Y(n21071) );
  XNOR2X1 U5717 ( .A(n3056), .B(n21058), .Y(n21072) );
  NOR2XL U5718 ( .A(n23884), .B(n26537), .Y(n4213) );
  CLKINVX3 U5719 ( .A(n22967), .Y(n3055) );
  CLKINVX8 U5720 ( .A(n3120), .Y(n3024) );
  CLKINVX3 U5721 ( .A(n22614), .Y(n3054) );
  INVX1 U5722 ( .A(n21852), .Y(n21265) );
  INVX2 U5723 ( .A(n3057), .Y(n3025) );
  BUFX16 U5724 ( .A(n11481), .Y(n21166) );
  CLKINVX3 U5725 ( .A(n22737), .Y(n3056) );
  OAI21X1 U5726 ( .A0(n14833), .A1(n26502), .B0(n14844), .Y(n14950) );
  CLKINVX3 U5727 ( .A(n22698), .Y(n3058) );
  NAND2X1 U5728 ( .A(n11172), .B(n11171), .Y(n22492) );
  NAND2X1 U5729 ( .A(n19346), .B(w2[31]), .Y(n8220) );
  AOI22X1 U5730 ( .A0(y11[23]), .A1(n19235), .B0(n19216), .B1(temp2[23]), .Y(
        n19214) );
  NAND2X1 U5731 ( .A(n19346), .B(w2[25]), .Y(n8083) );
  OAI21XL U5732 ( .A0(n26143), .A1(n21256), .B0(n21322), .Y(n21430) );
  AOI22X1 U5733 ( .A0(w2[93]), .A1(n19349), .B0(n3062), .B1(w1[125]), .Y(
        n14854) );
  AOI22X1 U5734 ( .A0(y11[26]), .A1(n19346), .B0(n3062), .B1(temp2[26]), .Y(
        n19229) );
  AOI22X1 U5735 ( .A0(n19346), .A1(w2[95]), .B0(n19216), .B1(w1[127]), .Y(
        n14963) );
  INVX1 U5736 ( .A(n22716), .Y(n22698) );
  NAND2X1 U5737 ( .A(n19346), .B(w2[30]), .Y(n7888) );
  INVX2 U5738 ( .A(n25059), .Y(n25820) );
  NAND2X1 U5739 ( .A(n19346), .B(w2[28]), .Y(n8101) );
  INVX8 U5740 ( .A(n3122), .Y(n3059) );
  CLKBUFX8 U5741 ( .A(n3063), .Y(n14833) );
  AOI22X1 U5742 ( .A0(y12[25]), .A1(n19346), .B0(n3026), .B1(temp3[25]), .Y(
        n14844) );
  NAND2X1 U5743 ( .A(n19346), .B(w2[29]), .Y(n8107) );
  NAND2X1 U5744 ( .A(n19346), .B(w2[26]), .Y(n8094) );
  AOI22X1 U5745 ( .A0(n19346), .A1(w2[63]), .B0(n3062), .B1(w1[95]), .Y(n19347) );
  NAND2X1 U5746 ( .A(n19346), .B(w2[27]), .Y(n8089) );
  INVX20 U5747 ( .A(n26595), .Y(n19346) );
  NAND2X1 U5748 ( .A(n11174), .B(n11173), .Y(n22491) );
  CLKINVX4 U5749 ( .A(n25428), .Y(n3064) );
  CLKINVX8 U5750 ( .A(n21111), .Y(n3026) );
  INVX8 U5751 ( .A(n26595), .Y(n3027) );
  CLKINVX4 U5752 ( .A(n4631), .Y(n21256) );
  INVX8 U5753 ( .A(n25428), .Y(n3028) );
  NAND2XL U5754 ( .A(in_valid_d), .B(w1[142]), .Y(n11530) );
  NOR2XL U5755 ( .A(n17167), .B(n25999), .Y(n5987) );
  INVXL U5756 ( .A(learning_rate[2]), .Y(n24000) );
  CLKINVX4 U5757 ( .A(valid[0]), .Y(n23973) );
  NAND2XL U5758 ( .A(in_valid_t), .B(learning_rate[25]), .Y(n11593) );
  CLKINVX3 U5759 ( .A(in_valid_w2), .Y(n23997) );
  INVX1 U5760 ( .A(data_point[2]), .Y(n6233) );
  INVX1 U5761 ( .A(n24864), .Y(n25407) );
  INVX1 U5762 ( .A(n24957), .Y(n25384) );
  INVX1 U5763 ( .A(n24909), .Y(n25392) );
  INVX1 U5764 ( .A(n24765), .Y(n25448) );
  INVX1 U5765 ( .A(n24839), .Y(n25421) );
  AOI2BB1XL U5766 ( .A0N(n25423), .A1N(n3118), .B0(n21016), .Y(n2217) );
  AOI2BB1XL U5767 ( .A0N(n25497), .A1N(n3118), .B0(n25043), .Y(n2211) );
  AOI2BB1XL U5768 ( .A0N(n25473), .A1N(n3118), .B0(n25045), .Y(n2213) );
  AOI2BB1XL U5769 ( .A0N(n25625), .A1N(n3118), .B0(n25033), .Y(n2201) );
  AOI2BB1XL U5770 ( .A0N(n25598), .A1N(n3118), .B0(n25035), .Y(n2203) );
  AOI2BB1XL U5771 ( .A0N(n25569), .A1N(n3118), .B0(n25037), .Y(n2205) );
  AOI2BB1XL U5772 ( .A0N(n25547), .A1N(n3118), .B0(n25039), .Y(n2207) );
  AOI22X1 U5773 ( .A0(n24692), .A1(n24860), .B0(n24908), .B1(n24816), .Y(
        n24817) );
  OAI2BB1XL U5774 ( .A0N(n20890), .A1N(n25385), .B0(n3601), .Y(n3600) );
  OAI2BB1XL U5775 ( .A0N(n20890), .A1N(n25393), .B0(n4814), .Y(n4813) );
  INVX1 U5776 ( .A(n24552), .Y(n25558) );
  AOI22XL U5777 ( .A0(n24692), .A1(n24725), .B0(n24908), .B1(n20264), .Y(
        n20265) );
  AOI2BB1XL U5778 ( .A0N(n25521), .A1N(n3118), .B0(n25041), .Y(n2209) );
  INVX1 U5779 ( .A(n24532), .Y(n25566) );
  AOI222XL U5780 ( .A0(n24644), .A1(n25744), .B0(n25743), .B1(y20[10]), .C0(
        n25509), .C1(n20890), .Y(n2370) );
  AOI22XL U5781 ( .A0(n24692), .A1(n24607), .B0(n24908), .B1(n24597), .Y(
        n24598) );
  XOR2X1 U5782 ( .A(n24883), .B(n24928), .Y(n24884) );
  AOI222XL U5783 ( .A0(n23701), .A1(n25744), .B0(n25743), .B1(y20[7]), .C0(
        n25546), .C1(n20890), .Y(n2367) );
  OAI21XL U5784 ( .A0(n25535), .A1(n3118), .B0(n25311), .Y(n2144) );
  AOI222XL U5785 ( .A0(n25740), .A1(n25744), .B0(n25743), .B1(y20[6]), .C0(
        n25739), .C1(n20890), .Y(n2366) );
  INVX1 U5786 ( .A(n24642), .Y(n25509) );
  INVX1 U5787 ( .A(n24741), .Y(n25460) );
  INVX1 U5788 ( .A(n25316), .Y(n25736) );
  INVX1 U5789 ( .A(n23656), .Y(n25496) );
  INVX1 U5790 ( .A(n25319), .Y(n25734) );
  XOR2X1 U5791 ( .A(n24586), .B(n24537), .Y(n24517) );
  XOR2X1 U5792 ( .A(n24495), .B(n24494), .Y(n24496) );
  NOR2X1 U5793 ( .A(n24953), .B(n24952), .Y(n25356) );
  XOR2X1 U5794 ( .A(n24562), .B(n23621), .Y(n20897) );
  NAND2X1 U5795 ( .A(n24531), .B(n20996), .Y(n24569) );
  NAND2X2 U5796 ( .A(n20379), .B(n20378), .Y(n20382) );
  INVX1 U5797 ( .A(n24956), .Y(n25353) );
  NAND2X1 U5798 ( .A(n24622), .B(n24618), .Y(n24658) );
  AOI21X1 U5799 ( .A0(n15928), .A1(n3077), .B0(n15896), .Y(n24591) );
  INVX1 U5800 ( .A(n4778), .Y(n4779) );
  NAND2X1 U5801 ( .A(n15900), .B(n3077), .Y(n21009) );
  AOI21X1 U5802 ( .A0(n24752), .A1(n3075), .B0(n20226), .Y(n24577) );
  NAND2X1 U5803 ( .A(n20864), .B(n23583), .Y(n20901) );
  NOR2X2 U5804 ( .A(n23226), .B(n22230), .Y(n23255) );
  INVX1 U5805 ( .A(n24793), .Y(n4778) );
  NOR2BX1 U5806 ( .AN(n15749), .B(n24400), .Y(n4443) );
  NAND2X1 U5807 ( .A(n20252), .B(n3075), .Y(n24856) );
  NAND2XL U5808 ( .A(n3069), .B(n20232), .Y(n20243) );
  NOR2X1 U5809 ( .A(n20560), .B(n8997), .Y(n20918) );
  XOR2X1 U5810 ( .A(n23339), .B(n23338), .Y(n23340) );
  XOR2X1 U5811 ( .A(n23314), .B(n23343), .Y(n23315) );
  OAI21XL U5812 ( .A0(n20574), .A1(n3073), .B0(n20573), .Y(n23833) );
  NOR2XL U5813 ( .A(n24399), .B(n15742), .Y(n15740) );
  OAI2BB1X1 U5814 ( .A0N(n20473), .A1N(n20501), .B0(n20500), .Y(n20537) );
  OAI22X1 U5815 ( .A0(n20202), .A1(n3072), .B0(n20149), .B1(n20138), .Y(n20230) );
  ADDFHX1 U5816 ( .A(n24291), .B(n3076), .CI(n15747), .CO(n15742), .S(n24292)
         );
  AOI21X1 U5817 ( .A0(n15839), .A1(n3070), .B0(n15768), .Y(n15858) );
  NAND2X1 U5818 ( .A(n15890), .B(n3077), .Y(n15815) );
  NOR2X1 U5819 ( .A(n15833), .B(n15832), .Y(n15866) );
  NOR2X1 U5820 ( .A(n20221), .B(n20220), .Y(n20239) );
  NOR2X1 U5821 ( .A(n20190), .B(n20189), .Y(n20248) );
  ADDFHX1 U5822 ( .A(n24073), .B(n3075), .CI(n20123), .CO(n20122), .S(n24068)
         );
  ADDFHX1 U5823 ( .A(n24058), .B(n3077), .CI(n15743), .CO(n15747), .S(n24059)
         );
  NOR2X1 U5824 ( .A(n15803), .B(n15802), .Y(n15843) );
  OAI21XL U5825 ( .A0(n25382), .A1(n3121), .B0(n20632), .Y(n2576) );
  AOI21XL U5826 ( .A0(n20489), .A1(n3071), .B0(n20393), .Y(n20506) );
  OAI22X1 U5827 ( .A0(n3127), .A1(n15807), .B0(n15760), .B1(n3070), .Y(n15882)
         );
  NAND2X2 U5828 ( .A(n22217), .B(n22212), .Y(n23224) );
  ADDFHX1 U5829 ( .A(n23859), .B(n3073), .CI(n8985), .CO(n8984), .S(n23857) );
  NAND2X1 U5830 ( .A(n9005), .B(n3071), .Y(n20508) );
  NOR2X1 U5831 ( .A(n20413), .B(n20412), .Y(n20482) );
  XOR2X1 U5832 ( .A(n23268), .B(n23267), .Y(n23269) );
  NOR2X1 U5833 ( .A(n20417), .B(n20416), .Y(n20484) );
  OAI21XL U5834 ( .A0(n22419), .A1(n22418), .B0(n22417), .Y(n23376) );
  AOI21X1 U5835 ( .A0(n22384), .A1(n3082), .B0(n22383), .Y(n23297) );
  ADDFHX1 U5836 ( .A(n23817), .B(n20576), .CI(n8986), .CO(n8985), .S(n23815)
         );
  OAI22XL U5837 ( .A0(n22270), .A1(n22269), .B0(n22461), .B1(n22268), .Y(
        n23341) );
  AOI21X1 U5838 ( .A0(n22414), .A1(n3082), .B0(n22369), .Y(n23318) );
  INVX8 U5839 ( .A(n24986), .Y(n3030) );
  NAND2X1 U5840 ( .A(n3067), .B(n9006), .Y(n9001) );
  NAND2X1 U5841 ( .A(n3067), .B(n9016), .Y(n8998) );
  NOR2BX1 U5842 ( .AN(n22172), .B(n22171), .Y(n22184) );
  ADDFHX1 U5843 ( .A(n23811), .B(n3068), .CI(n8987), .CO(n8986), .S(n23809) );
  AOI21X1 U5844 ( .A0(n25733), .A1(n3229), .B0(n4828), .Y(n23943) );
  NAND3BX1 U5845 ( .AN(n23392), .B(n22182), .C(n23232), .Y(n22183) );
  AOI21X1 U5846 ( .A0(n4456), .A1(n3135), .B0(n25270), .Y(n4455) );
  AOI2BB2XL U5847 ( .B0(n22176), .B1(n22175), .A0N(n22175), .A1N(n22176), .Y(
        n23392) );
  NAND2X1 U5848 ( .A(n22370), .B(n3079), .Y(n22381) );
  NAND2X1 U5849 ( .A(n22239), .B(n3082), .Y(n22268) );
  NAND2BXL U5850 ( .AN(n20826), .B(n4873), .Y(n4872) );
  NOR2X1 U5851 ( .A(n15761), .B(n3070), .Y(n15768) );
  OAI2BB1X1 U5852 ( .A0N(n19072), .A1N(n25807), .B0(n19071), .Y(n2614) );
  OAI21XL U5853 ( .A0(n4380), .A1(n3121), .B0(n4549), .Y(n2575) );
  NAND2BX1 U5854 ( .AN(n23910), .B(n23909), .Y(n23911) );
  NOR2X1 U5855 ( .A(n20298), .B(n20296), .Y(n20622) );
  NOR2X1 U5856 ( .A(n22308), .B(n23223), .Y(n22196) );
  CLKINVX3 U5857 ( .A(n20144), .Y(n20138) );
  AOI21X1 U5858 ( .A0(n8980), .A1(n8979), .B0(n8978), .Y(n8981) );
  OAI2BB1XL U5859 ( .A0N(n25807), .A1N(n3769), .B0(n20793), .Y(n2569) );
  CLKINVX3 U5860 ( .A(n15734), .Y(n25273) );
  NOR2X1 U5861 ( .A(n20822), .B(n20820), .Y(n23540) );
  INVX1 U5862 ( .A(n25483), .Y(n24673) );
  NAND2X1 U5863 ( .A(n24397), .B(n25767), .Y(n6021) );
  OAI21XL U5864 ( .A0(n24582), .A1(n4585), .B0(n4212), .Y(n2603) );
  NAND2XL U5865 ( .A(n3408), .B(n24245), .Y(n24246) );
  NAND2X1 U5866 ( .A(n4223), .B(n4221), .Y(n3860) );
  NOR2X1 U5867 ( .A(n20163), .B(n20162), .Y(n20164) );
  AOI2BB1X2 U5868 ( .A0N(n24147), .A1N(n3121), .B0(n4213), .Y(n4212) );
  AOI22XL U5869 ( .A0(n24277), .A1(n25807), .B0(n2984), .B1(temp2[27]), .Y(
        n24278) );
  BUFX3 U5870 ( .A(n23676), .Y(n25832) );
  AOI21XL U5871 ( .A0(n3882), .A1(n25767), .B0(n20320), .Y(n2266) );
  NOR2X1 U5872 ( .A(n24386), .B(n23664), .Y(n23665) );
  INVX1 U5873 ( .A(n24145), .Y(n24581) );
  NOR2X1 U5874 ( .A(n24386), .B(n24271), .Y(n24272) );
  NOR2X1 U5875 ( .A(n24386), .B(n24385), .Y(n24387) );
  NOR2X1 U5876 ( .A(n24228), .B(n25328), .Y(n24231) );
  NOR2XL U5877 ( .A(n24460), .B(n25255), .Y(n24257) );
  NOR2X1 U5878 ( .A(n24202), .B(n25328), .Y(n24205) );
  NAND2X1 U5879 ( .A(n3132), .B(n20991), .Y(n20992) );
  BUFX12 U5880 ( .A(n23883), .Y(n3081) );
  MXI2X1 U5881 ( .A(n24249), .B(n20940), .S0(n4875), .Y(n20941) );
  INVXL U5882 ( .A(n25007), .Y(n3135) );
  AOI31X1 U5883 ( .A0(n22161), .A1(n22140), .A2(n22164), .B0(n22139), .Y(
        n22281) );
  NAND2X1 U5884 ( .A(n4219), .B(n3858), .Y(n4218) );
  NAND2X1 U5885 ( .A(n23808), .B(n5559), .Y(n3550) );
  MXI2XL U5886 ( .A(mul5_out[24]), .B(n25200), .S0(n3111), .Y(n2344) );
  MXI2XL U5887 ( .A(mul5_out[25]), .B(n25192), .S0(n3111), .Y(n2346) );
  INVX2 U5888 ( .A(n23509), .Y(n23579) );
  OR2X2 U5889 ( .A(n15801), .B(n15809), .Y(n15722) );
  INVX1 U5890 ( .A(n3014), .Y(n4219) );
  AOI2BB1XL U5891 ( .A0N(n22146), .A1N(n22273), .B0(n22272), .Y(n22147) );
  NAND2XL U5892 ( .A(n17436), .B(n5720), .Y(n5701) );
  XOR2X1 U5893 ( .A(n15673), .B(n15672), .Y(n15801) );
  OAI21XL U5894 ( .A0(n25222), .A1(n23636), .B0(n25221), .Y(mul5_out[23]) );
  NAND3X1 U5895 ( .A(n23734), .B(n4185), .C(n18972), .Y(n23735) );
  NOR3X2 U5896 ( .A(n3318), .B(n3320), .C(n3308), .Y(n3235) );
  NAND2XL U5897 ( .A(n23514), .B(n23734), .Y(n23517) );
  NAND2X1 U5898 ( .A(n4508), .B(n4651), .Y(n23565) );
  INVX1 U5899 ( .A(n25294), .Y(n25330) );
  NOR2XL U5900 ( .A(n23573), .B(n23572), .Y(n3667) );
  NAND3X2 U5901 ( .A(n4648), .B(n20714), .C(n20614), .Y(n3321) );
  NAND2X1 U5902 ( .A(n8651), .B(n8918), .Y(n8653) );
  XOR2X1 U5903 ( .A(n5573), .B(n20619), .Y(n23806) );
  AOI21X1 U5904 ( .A0(n8635), .A1(n8889), .B0(n8634), .Y(n8758) );
  NAND2X1 U5905 ( .A(n3895), .B(n20323), .Y(n20325) );
  INVX1 U5906 ( .A(n20715), .Y(n5524) );
  INVXL U5907 ( .A(n15640), .Y(n15655) );
  INVX1 U5908 ( .A(n4305), .Y(n20270) );
  XOR2X1 U5909 ( .A(n20361), .B(n20360), .Y(n20942) );
  INVX1 U5910 ( .A(n8905), .Y(n8941) );
  BUFX8 U5911 ( .A(n3938), .Y(n3895) );
  NAND2X1 U5912 ( .A(n19779), .B(n20047), .Y(n19781) );
  INVX1 U5913 ( .A(n20617), .Y(n5600) );
  XOR2X1 U5914 ( .A(n20746), .B(n20745), .Y(n21052) );
  NAND2X1 U5915 ( .A(n15398), .B(n15668), .Y(n15400) );
  OAI21X1 U5916 ( .A0(n15372), .A1(n15656), .B0(n15371), .Y(n15640) );
  XNOR2X1 U5917 ( .A(n20071), .B(n20070), .Y(n20156) );
  NOR2XL U5918 ( .A(n20929), .B(n20928), .Y(n20930) );
  NAND2XL U5919 ( .A(n3357), .B(n20359), .Y(n20361) );
  NAND3X2 U5920 ( .A(n3339), .B(n3337), .C(n3336), .Y(n3806) );
  CLKINVX2 U5921 ( .A(n17434), .Y(n17437) );
  NAND2X1 U5922 ( .A(n5100), .B(n20868), .Y(n20871) );
  INVX1 U5923 ( .A(n8927), .Y(n8912) );
  NOR2XL U5924 ( .A(n9000), .B(n8999), .Y(n8943) );
  AND2X1 U5925 ( .A(n23486), .B(n6222), .Y(n25335) );
  NAND2X1 U5926 ( .A(n3596), .B(n5100), .Y(n20758) );
  NOR2XL U5927 ( .A(n15642), .B(n15643), .Y(n15382) );
  NAND4X2 U5928 ( .A(n4416), .B(n4652), .C(n4994), .D(n23749), .Y(n3379) );
  NAND4X2 U5929 ( .A(n4076), .B(n13037), .C(n13024), .D(n20671), .Y(n4414) );
  NAND2X1 U5930 ( .A(n20857), .B(n5100), .Y(n20859) );
  AOI21X1 U5931 ( .A0(n15208), .A1(n15378), .B0(n15377), .Y(n15641) );
  XOR2X1 U5932 ( .A(n19078), .B(n19077), .Y(n20907) );
  INVXL U5933 ( .A(n13037), .Y(n4060) );
  INVX1 U5934 ( .A(n23529), .Y(n23530) );
  INVX1 U5935 ( .A(n3958), .Y(n20927) );
  AOI21X1 U5936 ( .A0(n19738), .A1(n19759), .B0(n19758), .Y(n20019) );
  NAND2XL U5937 ( .A(n20920), .B(n5394), .Y(n17468) );
  NAND2XL U5938 ( .A(n15695), .B(n15694), .Y(n15656) );
  NAND2XL U5939 ( .A(n20074), .B(n20072), .Y(n20034) );
  CLKINVX3 U5940 ( .A(n2999), .Y(n3144) );
  INVX1 U5941 ( .A(n10597), .Y(n10598) );
  NAND2X1 U5942 ( .A(n15662), .B(n15682), .Y(n15392) );
  INVX1 U5943 ( .A(n18830), .Y(n6033) );
  INVX1 U5944 ( .A(n21947), .Y(n22117) );
  NAND4BX2 U5945 ( .AN(n20312), .B(n3145), .C(n13028), .D(n13026), .Y(n4413)
         );
  BUFX8 U5946 ( .A(n3848), .Y(n3357) );
  AOI21X1 U5947 ( .A0(n22077), .A1(n21820), .B0(n21819), .Y(n21947) );
  NOR2XL U5948 ( .A(n21039), .B(n5410), .Y(n3668) );
  NAND2X1 U5949 ( .A(n15384), .B(n15383), .Y(n15676) );
  INVX1 U5950 ( .A(n10972), .Y(n10982) );
  INVX1 U5951 ( .A(n15677), .Y(n15662) );
  OR2X2 U5952 ( .A(n8641), .B(n8640), .Y(n8403) );
  CLKINVX3 U5953 ( .A(n21039), .Y(n3145) );
  NAND2X2 U5954 ( .A(n23454), .B(n6024), .Y(n23476) );
  INVX1 U5955 ( .A(n20056), .Y(n20041) );
  NOR2X1 U5956 ( .A(n20141), .B(n20147), .Y(n20074) );
  NAND2BX1 U5957 ( .AN(n8622), .B(n4815), .Y(n8908) );
  NAND2X1 U5958 ( .A(n19765), .B(n19764), .Y(n20055) );
  NAND2X1 U5959 ( .A(n6030), .B(n4675), .Y(n6029) );
  NAND2X2 U5960 ( .A(n20348), .B(n20926), .Y(n3329) );
  NAND4X2 U5961 ( .A(n3010), .B(n17466), .C(n17421), .D(n17455), .Y(n3931) );
  INVX1 U5962 ( .A(n15589), .Y(n15628) );
  INVX1 U5963 ( .A(n20279), .Y(n20856) );
  INVXL U5964 ( .A(n17471), .Y(n5711) );
  NAND2X1 U5965 ( .A(n8813), .B(n8812), .Y(n8843) );
  OR2X2 U5966 ( .A(n15388), .B(n15387), .Y(n15682) );
  NAND2X1 U5967 ( .A(n10635), .B(n10574), .Y(n3317) );
  NOR2XL U5968 ( .A(n20891), .B(n20896), .Y(n20892) );
  INVX1 U5969 ( .A(n10627), .Y(n10628) );
  OR2XL U5970 ( .A(n20952), .B(n20951), .Y(n20953) );
  NAND2X1 U5971 ( .A(n20145), .B(n19952), .Y(n20147) );
  NOR2BXL U5972 ( .AN(n5220), .B(n10608), .Y(n4072) );
  NAND2X2 U5973 ( .A(n20894), .B(n3536), .Y(n20279) );
  NOR2X1 U5974 ( .A(n15565), .B(n15564), .Y(n15589) );
  AND2X4 U5975 ( .A(n17466), .B(n17435), .Y(n3956) );
  OAI2BB1XL U5976 ( .A0N(n18917), .A1N(n18918), .B0(n4507), .Y(n4407) );
  OAI21XL U5977 ( .A0(n8600), .A1(n8599), .B0(n8598), .Y(n9004) );
  OR2X2 U5978 ( .A(n19769), .B(n19768), .Y(n19534) );
  NAND2X1 U5979 ( .A(n15567), .B(n15566), .Y(n15634) );
  OR2X1 U5980 ( .A(n8417), .B(n8614), .Y(n8419) );
  INVX1 U5981 ( .A(n3748), .Y(n13030) );
  XOR2X1 U5982 ( .A(n4623), .B(n22186), .Y(n22198) );
  OR2X1 U5983 ( .A(n8614), .B(n8440), .Y(n8442) );
  INVX1 U5984 ( .A(n20762), .Y(n20763) );
  NOR2X2 U5985 ( .A(n12908), .B(n12929), .Y(n4411) );
  NOR2X2 U5986 ( .A(n12904), .B(n12929), .Y(n3349) );
  NAND3X1 U5987 ( .A(n10741), .B(n10739), .C(n20277), .Y(n3526) );
  INVX1 U5988 ( .A(n19968), .Y(n20007) );
  NAND2X1 U5989 ( .A(n22099), .B(n6202), .Y(n21830) );
  NOR2X1 U5990 ( .A(n19944), .B(n19943), .Y(n19968) );
  NAND2X1 U5991 ( .A(n19946), .B(n19945), .Y(n20013) );
  NAND2X1 U5992 ( .A(n4051), .B(n12809), .Y(n12818) );
  NAND2X2 U5993 ( .A(n18792), .B(n3007), .Y(n3355) );
  INVXL U5994 ( .A(n20744), .Y(n20745) );
  OR2X1 U5995 ( .A(n15359), .B(n15123), .Y(n15125) );
  OAI2BB1XL U5996 ( .A0N(n12892), .A1N(n12914), .B0(n12891), .Y(n12894) );
  OR2XL U5997 ( .A(n19595), .B(n19748), .Y(n19597) );
  OR2X1 U5998 ( .A(n19748), .B(n19505), .Y(n19507) );
  NAND2X1 U5999 ( .A(n17356), .B(n17355), .Y(n3809) );
  INVX1 U6000 ( .A(n20277), .Y(n20880) );
  NAND2BXL U6001 ( .AN(n12928), .B(n12892), .Y(n4012) );
  INVX1 U6002 ( .A(n10739), .Y(n20275) );
  NOR2X2 U6003 ( .A(n10603), .B(n10479), .Y(n10480) );
  NAND2X1 U6004 ( .A(n4131), .B(n17329), .Y(n4130) );
  NAND2X1 U6005 ( .A(n8295), .B(n8790), .Y(n8792) );
  AOI21X1 U6006 ( .A0(n8807), .A1(n8823), .B0(n3155), .Y(n8806) );
  NOR4BXL U6007 ( .AN(n15344), .B(n15343), .C(n15342), .D(n15341), .Y(n15346)
         );
  INVX1 U6008 ( .A(n11393), .Y(n11372) );
  AOI21X1 U6009 ( .A0(n21967), .A1(n22042), .B0(n21966), .Y(n21968) );
  OAI21XL U6010 ( .A0(n19685), .A1(n19684), .B0(n19683), .Y(n19686) );
  XOR2X2 U6011 ( .A(n7326), .B(n3566), .Y(n20896) );
  INVX1 U6012 ( .A(n3781), .Y(n3688) );
  NAND2BX1 U6013 ( .AN(n17337), .B(n3781), .Y(n3334) );
  AOI2BB1X2 U6014 ( .A0N(n17306), .A1N(n17305), .B0(n4149), .Y(n3959) );
  CLKINVX3 U6015 ( .A(n17419), .Y(n3085) );
  NAND2X1 U6016 ( .A(n15046), .B(n15549), .Y(n15551) );
  NAND2X1 U6017 ( .A(n12864), .B(n12827), .Y(n12828) );
  NAND2X1 U6018 ( .A(n15046), .B(n15544), .Y(n15546) );
  CLKINVX3 U6019 ( .A(n3781), .Y(n3335) );
  NAND2X1 U6020 ( .A(n14592), .B(n14591), .Y(n14593) );
  NAND2XL U6021 ( .A(n12845), .B(n12840), .Y(n4917) );
  XNOR2X1 U6022 ( .A(n7007), .B(n7006), .Y(n10738) );
  NAND2X1 U6023 ( .A(n20641), .B(n20642), .Y(n20643) );
  NAND2X1 U6024 ( .A(n14626), .B(n14625), .Y(n14627) );
  AND2X2 U6025 ( .A(n10221), .B(n10220), .Y(n4613) );
  AOI2BB2XL U6026 ( .B0(n8435), .B1(n3157), .A0N(n3157), .A1N(n8431), .Y(n8517) );
  NAND2X1 U6027 ( .A(n5667), .B(n17370), .Y(n5059) );
  AOI2BB2XL U6028 ( .B0(n3087), .B1(n8435), .A0N(n8434), .A1N(n8433), .Y(n8655) );
  AND2X2 U6029 ( .A(n10188), .B(n10187), .Y(n4614) );
  AND2X2 U6030 ( .A(n18921), .B(n18920), .Y(n18922) );
  NOR2X1 U6031 ( .A(n15350), .B(n3090), .Y(n15572) );
  INVX1 U6032 ( .A(n14603), .Y(n14626) );
  NOR2X1 U6033 ( .A(n19592), .B(n19807), .Y(n19898) );
  AND2X2 U6034 ( .A(n10245), .B(n10244), .Y(n4603) );
  AND2X1 U6035 ( .A(n15424), .B(n15336), .Y(n15549) );
  NOR2X1 U6036 ( .A(n15408), .B(n3090), .Y(n15539) );
  AOI2BB2X1 U6037 ( .B0(n19475), .B1(n19542), .A0N(n19542), .A1N(n19536), .Y(
        n19592) );
  INVX1 U6038 ( .A(n10208), .Y(n10245) );
  NOR2X1 U6039 ( .A(n21887), .B(n21886), .Y(n21921) );
  INVXL U6040 ( .A(n10466), .Y(n4360) );
  NAND2X1 U6041 ( .A(n22004), .B(n22003), .Y(n22064) );
  NOR2X1 U6042 ( .A(n22004), .B(n22003), .Y(n22027) );
  NAND2X1 U6043 ( .A(n10227), .B(n10230), .Y(n4640) );
  AOI2BB2XL U6044 ( .B0(n3087), .B1(n8412), .A0N(n3087), .A1N(n8404), .Y(n8502) );
  NAND2X1 U6045 ( .A(n13999), .B(n13998), .Y(n14586) );
  INVX1 U6046 ( .A(n9197), .Y(n9198) );
  NAND2BX1 U6047 ( .AN(n8555), .B(n8592), .Y(n8603) );
  NAND2X1 U6048 ( .A(n12978), .B(n12858), .Y(n12861) );
  OR2X1 U6049 ( .A(n21597), .B(n21787), .Y(n21599) );
  NAND2XL U6050 ( .A(n3157), .B(n8571), .Y(n8551) );
  ADDFHX1 U6051 ( .A(n10445), .B(n10444), .CI(n10443), .CO(n10468), .S(n10466)
         );
  NAND2X1 U6052 ( .A(n14564), .B(n14563), .Y(n14565) );
  CLKINVX3 U6053 ( .A(n19807), .Y(n3159) );
  AND2X2 U6054 ( .A(n14654), .B(n14659), .Y(n4636) );
  INVX1 U6055 ( .A(n7823), .Y(n7824) );
  INVX4 U6056 ( .A(n8434), .Y(n3157) );
  OAI21X1 U6057 ( .A0(n4232), .A1(n4229), .B0(n4228), .Y(n5367) );
  CLKINVX3 U6058 ( .A(n14313), .Y(n3088) );
  INVX1 U6059 ( .A(n3422), .Y(n17214) );
  OR2X2 U6060 ( .A(n17320), .B(n4104), .Y(n4102) );
  INVX1 U6061 ( .A(n17252), .Y(n17254) );
  AOI21X1 U6062 ( .A0(n21996), .A1(n3222), .B0(n21849), .Y(n21995) );
  INVX1 U6063 ( .A(n15277), .Y(n15303) );
  NAND2XL U6064 ( .A(n3278), .B(n3277), .Y(n3276) );
  NAND2X1 U6065 ( .A(n14543), .B(n14541), .Y(n14530) );
  AND2X2 U6066 ( .A(n10625), .B(n10624), .Y(n4607) );
  NAND2X2 U6067 ( .A(n3720), .B(n12873), .Y(n3719) );
  INVXL U6068 ( .A(n4676), .Y(n3274) );
  XOR2X1 U6069 ( .A(n6165), .B(n10429), .Y(n10319) );
  AOI21X1 U6070 ( .A0(n18928), .A1(n18932), .B0(n18935), .Y(n18929) );
  INVX2 U6071 ( .A(n3090), .Y(n3034) );
  AOI21X1 U6072 ( .A0(n13034), .A1(n13033), .B0(n13032), .Y(n13035) );
  INVX1 U6073 ( .A(n7013), .Y(n7015) );
  AND2X2 U6074 ( .A(n12893), .B(n12907), .Y(n4629) );
  CLKINVX3 U6075 ( .A(n14314), .Y(n3089) );
  NAND2X1 U6076 ( .A(n12862), .B(n12863), .Y(n4612) );
  NAND2X1 U6077 ( .A(n5379), .B(n10083), .Y(n5378) );
  NAND2X1 U6078 ( .A(n21506), .B(n21989), .Y(n21991) );
  NAND2X1 U6079 ( .A(n12837), .B(n12779), .Y(n4037) );
  INVXL U6080 ( .A(n4304), .Y(n4175) );
  AND2X2 U6081 ( .A(n4943), .B(n17314), .Y(n4646) );
  NAND2BX1 U6082 ( .AN(n19644), .B(n3094), .Y(n19688) );
  NAND2X1 U6083 ( .A(n10474), .B(n10473), .Y(n10630) );
  ADDFHX1 U6084 ( .A(n9485), .B(n9484), .CI(n9483), .CO(n9489), .S(n9486) );
  NAND2XL U6085 ( .A(n10555), .B(n10645), .Y(n4676) );
  OAI21X1 U6086 ( .A0(n7822), .A1(n7821), .B0(n7820), .Y(n7823) );
  NAND2XL U6087 ( .A(n3280), .B(n9764), .Y(n3275) );
  AOI21X1 U6088 ( .A0(n18928), .A1(n18847), .B0(n18851), .Y(n18852) );
  AOI2BB2XL U6089 ( .B0(n21864), .B1(n3096), .A0N(n3096), .A1N(n21603), .Y(
        n21641) );
  AND2X2 U6090 ( .A(n10601), .B(n10600), .Y(n4687) );
  NAND2X2 U6091 ( .A(n17122), .B(n17339), .Y(n4104) );
  AOI21X1 U6092 ( .A0(n18981), .A1(n18709), .B0(n18708), .Y(n19008) );
  OAI21XL U6093 ( .A0(n8252), .A1(n8267), .B0(n8269), .Y(n8227) );
  NAND2X1 U6094 ( .A(n4949), .B(n12915), .Y(n4594) );
  INVX1 U6095 ( .A(n7321), .Y(n7322) );
  AOI2BB2X1 U6096 ( .B0(n21783), .B1(n3096), .A0N(n3096), .A1N(n21782), .Y(
        n21846) );
  AOI21X1 U6097 ( .A0(n7321), .A1(n7325), .B0(n7309), .Y(n7310) );
  NAND2XL U6098 ( .A(n5390), .B(n4323), .Y(n9483) );
  INVXL U6099 ( .A(n7019), .Y(n7009) );
  INVXL U6100 ( .A(n7018), .Y(n7010) );
  ADDFHX1 U6101 ( .A(n10442), .B(n10441), .CI(n10440), .CO(n10472), .S(n10469)
         );
  ADDFHX2 U6102 ( .A(n16784), .B(n16782), .CI(n16783), .CO(n16850), .S(n16849)
         );
  NAND2X1 U6103 ( .A(n12111), .B(n3472), .Y(n3471) );
  NAND2X1 U6104 ( .A(n15025), .B(n15024), .Y(n15029) );
  INVXL U6105 ( .A(n17372), .Y(n17373) );
  INVXL U6106 ( .A(n14484), .Y(n14539) );
  NAND2X1 U6107 ( .A(n14516), .B(n14515), .Y(n14517) );
  AOI2BB2XL U6108 ( .B0(n21571), .B1(n3096), .A0N(n3096), .A1N(n21766), .Y(
        n21659) );
  AOI21X1 U6109 ( .A0(n11000), .A1(n10950), .B0(n10949), .Y(n11021) );
  AND2X2 U6110 ( .A(n18947), .B(n18945), .Y(n4593) );
  OR2X2 U6111 ( .A(n10052), .B(n10051), .Y(n9762) );
  INVX1 U6112 ( .A(n7236), .Y(n5622) );
  XOR2X1 U6113 ( .A(n4459), .B(n4458), .Y(n4457) );
  NAND2XL U6114 ( .A(n10317), .B(n10318), .Y(n5221) );
  OR2X2 U6115 ( .A(n12773), .B(n12772), .Y(n12611) );
  INVX1 U6116 ( .A(n10439), .Y(n3163) );
  NAND2XL U6117 ( .A(n3096), .B(n21696), .Y(n21707) );
  NAND2XL U6118 ( .A(n9716), .B(n9717), .Y(n5140) );
  OAI21X1 U6119 ( .A0(n6100), .A1(n6099), .B0(n6097), .Y(n14067) );
  AND2X2 U6120 ( .A(n7426), .B(n7424), .Y(n7318) );
  NOR2X1 U6121 ( .A(n14328), .B(n14327), .Y(n14484) );
  INVXL U6122 ( .A(n4316), .Y(n4315) );
  NAND2X1 U6123 ( .A(n14272), .B(n14495), .Y(n14335) );
  NAND2X1 U6124 ( .A(n14272), .B(n14499), .Y(n14500) );
  ADDFHX1 U6125 ( .A(n17958), .B(n17957), .CI(n17956), .CO(n18321), .S(n18320)
         );
  NAND2X1 U6126 ( .A(n17113), .B(n17112), .Y(n17332) );
  INVX1 U6127 ( .A(n17338), .Y(n17321) );
  AOI22X1 U6128 ( .A0(n3095), .A1(n21592), .B0(n21643), .B1(n21580), .Y(n21864) );
  CLKINVX3 U6129 ( .A(n3096), .Y(n3172) );
  NAND2X1 U6130 ( .A(n18686), .B(n18685), .Y(n18945) );
  NAND2X1 U6131 ( .A(n17118), .B(n17117), .Y(n17342) );
  NAND2X1 U6132 ( .A(n17115), .B(n17116), .Y(n17338) );
  NOR2X2 U6133 ( .A(n17118), .B(n17117), .Y(n17326) );
  NAND2X2 U6134 ( .A(n6908), .B(n6907), .Y(n7366) );
  INVX1 U6135 ( .A(n7317), .Y(n7426) );
  NAND2X1 U6136 ( .A(n3897), .B(n3899), .Y(n3896) );
  INVX1 U6137 ( .A(n16780), .Y(n3611) );
  NOR2X1 U6138 ( .A(n12866), .B(n12788), .Y(n12807) );
  OAI21XL U6139 ( .A0(n5040), .A1(n5039), .B0(n5038), .Y(n12773) );
  XNOR3X2 U6140 ( .A(n3474), .B(n12112), .C(n12111), .Y(n12424) );
  OR2XL U6141 ( .A(n10005), .B(n10004), .Y(n10003) );
  NAND2X1 U6142 ( .A(n3902), .B(n3898), .Y(n3897) );
  NAND2X1 U6143 ( .A(n17120), .B(n17119), .Y(n17349) );
  OAI21X2 U6144 ( .A0(n5831), .A1(n5830), .B0(n5829), .Y(n17118) );
  OAI2BB1X1 U6145 ( .A0N(n17004), .A1N(n17003), .B0(n4100), .Y(n17012) );
  XNOR2X1 U6146 ( .A(n16954), .B(n5687), .Y(n17115) );
  ADDFHX1 U6147 ( .A(n9805), .B(n9804), .CI(n9803), .CO(n9830), .S(n9806) );
  NAND2XL U6148 ( .A(n12688), .B(n12689), .Y(n6113) );
  NAND2X1 U6149 ( .A(n19406), .B(n19405), .Y(n19407) );
  NAND2X2 U6150 ( .A(n3799), .B(n3798), .Y(n16224) );
  INVXL U6151 ( .A(n12976), .Y(n12868) );
  XOR2X2 U6152 ( .A(n3742), .B(n12475), .Y(n12484) );
  OAI21X1 U6153 ( .A0(n12480), .A1(n12481), .B0(n3908), .Y(n3905) );
  NAND2X1 U6154 ( .A(n12775), .B(n12774), .Y(n12849) );
  NAND2XL U6155 ( .A(n5350), .B(n5349), .Y(n9294) );
  NAND2X1 U6156 ( .A(n5774), .B(n5773), .Y(n11858) );
  ADDFHX2 U6157 ( .A(n10294), .B(n10293), .CI(n10292), .CO(n10430), .S(n10316)
         );
  NAND2X1 U6158 ( .A(n7484), .B(n7488), .Y(n7485) );
  NAND3BXL U6159 ( .AN(n6665), .B(n6658), .C(n4635), .Y(n5556) );
  NAND2XL U6160 ( .A(n6893), .B(n5613), .Y(n5612) );
  NOR2X1 U6161 ( .A(M6_mult_x_15_n462), .B(M6_mult_x_15_n457), .Y(n10973) );
  OR2X2 U6162 ( .A(n14343), .B(n14342), .Y(n14651) );
  OR2X1 U6163 ( .A(M6_mult_x_15_n469), .B(M6_mult_x_15_n475), .Y(n11000) );
  NAND2X1 U6164 ( .A(n23844), .B(n8281), .Y(n8285) );
  NOR2X1 U6165 ( .A(n23158), .B(n23157), .Y(n14960) );
  NAND2BX1 U6166 ( .AN(n10721), .B(n7420), .Y(n7872) );
  INVX1 U6167 ( .A(n7877), .Y(n7873) );
  OAI21X1 U6168 ( .A0(n16169), .A1(n16170), .B0(n3800), .Y(n3799) );
  XOR2X2 U6169 ( .A(n16805), .B(n16804), .Y(n3421) );
  INVX1 U6170 ( .A(n5396), .Y(n7764) );
  AND2X2 U6171 ( .A(n6729), .B(n6730), .Y(n3480) );
  INVX1 U6172 ( .A(n23182), .Y(n8224) );
  XNOR2X1 U6173 ( .A(n21468), .B(n21467), .Y(n21560) );
  AOI21X1 U6174 ( .A0(n7806), .A1(n7812), .B0(n7679), .Y(n7680) );
  INVXL U6175 ( .A(n16804), .Y(n3683) );
  NAND2X1 U6176 ( .A(n12683), .B(n12682), .Y(n5929) );
  NOR2XL U6177 ( .A(n24045), .B(n24044), .Y(n4499) );
  OAI21X2 U6178 ( .A0(n3343), .A1(n3342), .B0(n3341), .Y(n16138) );
  INVX1 U6179 ( .A(n7657), .Y(n7771) );
  ADDFHX1 U6180 ( .A(n17022), .B(n17021), .CI(n17020), .CO(n17029), .S(n17027)
         );
  ADDFHX1 U6181 ( .A(n17010), .B(n17009), .CI(n17008), .CO(n17116), .S(n17113)
         );
  NAND2BXL U6182 ( .AN(n6894), .B(n5614), .Y(n5613) );
  INVX1 U6183 ( .A(n6119), .Y(n3340) );
  NAND2X1 U6184 ( .A(n23642), .B(n23641), .Y(n23644) );
  INVXL U6185 ( .A(n16767), .Y(n3942) );
  CLKINVX8 U6186 ( .A(n3094), .Y(n3039) );
  INVX1 U6187 ( .A(n12480), .Y(n3906) );
  OAI21X2 U6188 ( .A0(n3651), .A1(n4133), .B0(n3650), .Y(n3908) );
  INVX1 U6189 ( .A(n11824), .Y(n4025) );
  ADDFHX1 U6190 ( .A(n11828), .B(n11827), .CI(n11826), .CO(n11823), .S(n12474)
         );
  INVX1 U6191 ( .A(n18315), .Y(n3097) );
  INVX1 U6192 ( .A(n18980), .Y(n19004) );
  NAND2X1 U6193 ( .A(M6_mult_x_15_n445), .B(M6_mult_x_15_n442), .Y(n11008) );
  ADDFHX2 U6194 ( .A(n17726), .B(n17725), .CI(n17724), .CO(n17688), .S(n18332)
         );
  NAND2XL U6195 ( .A(n12376), .B(n12383), .Y(n4237) );
  ADDFHX1 U6196 ( .A(n9476), .B(n9475), .CI(n9474), .CO(n9522), .S(n9453) );
  ADDFHX1 U6197 ( .A(n10079), .B(n10078), .CI(n10077), .CO(n10103), .S(n10093)
         );
  ADDFHX2 U6198 ( .A(n12465), .B(n12464), .CI(n12463), .CO(n12486), .S(n12466)
         );
  AND2X2 U6199 ( .A(n7786), .B(n7785), .Y(n4641) );
  NAND2X1 U6200 ( .A(n12784), .B(n12783), .Y(n12976) );
  INVXL U6201 ( .A(n14022), .Y(n6100) );
  NOR2XL U6202 ( .A(n12676), .B(n12677), .Y(n3980) );
  OR2X1 U6203 ( .A(M6_mult_x_15_n434), .B(n11093), .Y(n11367) );
  OAI21XL U6204 ( .A0(n11720), .A1(n11719), .B0(n11718), .Y(n4427) );
  INVXL U6205 ( .A(n11720), .Y(n4429) );
  OAI2BB1X1 U6206 ( .A0N(n4317), .A1N(n4509), .B0(n17595), .Y(n3428) );
  XOR3X2 U6207 ( .A(n11791), .B(n11790), .C(n11789), .Y(n11866) );
  NAND2X1 U6208 ( .A(n4958), .B(n4957), .Y(n11768) );
  INVXL U6209 ( .A(n4509), .Y(n4183) );
  ADDFHX2 U6210 ( .A(n11838), .B(n11837), .CI(n11836), .CO(n11826), .S(n12480)
         );
  NAND2XL U6211 ( .A(n6079), .B(n17550), .Y(n6078) );
  NAND2X1 U6212 ( .A(n7703), .B(n7724), .Y(n7699) );
  ADDFHX2 U6213 ( .A(n17955), .B(n17954), .CI(n17953), .CO(n18384), .S(n17956)
         );
  XOR2X2 U6214 ( .A(n16434), .B(n16433), .Y(n3706) );
  NAND2X1 U6215 ( .A(n17126), .B(n17125), .Y(n17351) );
  AND2X2 U6216 ( .A(n7812), .B(n7811), .Y(n4691) );
  XNOR3X2 U6217 ( .A(n17596), .B(n4509), .C(n17595), .Y(n17692) );
  NAND2XL U6218 ( .A(n17918), .B(n5813), .Y(n4069) );
  NAND2X1 U6219 ( .A(n16300), .B(n16301), .Y(n5330) );
  INVX1 U6220 ( .A(n3955), .Y(n3954) );
  AND2XL U6221 ( .A(n6669), .B(n6668), .Y(n6670) );
  INVX1 U6222 ( .A(n23161), .Y(n14970) );
  INVX1 U6223 ( .A(n23162), .Y(n14969) );
  INVX1 U6224 ( .A(n23163), .Y(n14968) );
  INVX1 U6225 ( .A(n23164), .Y(n14979) );
  XNOR2X1 U6226 ( .A(n11920), .B(n4974), .Y(n3658) );
  INVX1 U6227 ( .A(n23160), .Y(n15017) );
  ADDFHX2 U6228 ( .A(n6809), .B(n6808), .CI(n6807), .CO(n6903), .S(n6810) );
  NAND2X1 U6229 ( .A(n18705), .B(n18704), .Y(n19003) );
  NAND2XL U6230 ( .A(n16762), .B(n16763), .Y(n3946) );
  INVX1 U6231 ( .A(n12812), .Y(n12817) );
  AOI22XL U6232 ( .A0(n18267), .A1(n18266), .B0(n18264), .B1(n18265), .Y(
        n18268) );
  NAND2XL U6233 ( .A(n9377), .B(n3266), .Y(n3265) );
  NAND2X1 U6234 ( .A(n4020), .B(n6003), .Y(n4019) );
  NAND2X1 U6235 ( .A(n7664), .B(n7663), .Y(n7762) );
  NAND2X1 U6236 ( .A(n21447), .B(n21479), .Y(n21448) );
  AOI21X1 U6237 ( .A0(n21484), .A1(n21483), .B0(n21482), .Y(n21505) );
  NAND2XL U6238 ( .A(n3822), .B(n3821), .Y(n17800) );
  INVX1 U6239 ( .A(n7749), .Y(n7806) );
  ADDFHX2 U6240 ( .A(n12462), .B(n12461), .CI(n12460), .CO(n12467), .S(n12469)
         );
  INVX1 U6241 ( .A(n21483), .Y(n21468) );
  ADDFHX1 U6242 ( .A(n18101), .B(n18099), .CI(n18100), .CO(n18306), .S(n18302)
         );
  NAND2XL U6243 ( .A(n12134), .B(n3385), .Y(n3384) );
  OAI21X1 U6244 ( .A0(n14120), .A1(n13861), .B0(n5487), .Y(n13849) );
  NAND2XL U6245 ( .A(n5369), .B(n5368), .Y(n12650) );
  NAND2BXL U6246 ( .AN(n10157), .B(n3099), .Y(n4358) );
  OAI22XL U6247 ( .A0(n15548), .A1(n3101), .B0(n15558), .B1(n15547), .Y(n15564) );
  NAND2BXL U6248 ( .AN(n9208), .B(n3099), .Y(n4339) );
  NAND2BXL U6249 ( .AN(n9653), .B(n3099), .Y(n5149) );
  CLKINVX2 U6250 ( .A(n16171), .Y(n3369) );
  ADDFHX2 U6251 ( .A(n6416), .B(n6415), .CI(n6414), .CO(n6388), .S(n6418) );
  NAND2X1 U6252 ( .A(n11692), .B(n4959), .Y(n4958) );
  NAND2BX1 U6253 ( .AN(n10367), .B(n3297), .Y(n3296) );
  INVX1 U6254 ( .A(n23209), .Y(n19352) );
  INVX1 U6255 ( .A(n23206), .Y(n19403) );
  INVX1 U6256 ( .A(n23208), .Y(n19353) );
  NAND2X1 U6257 ( .A(n8482), .B(n8184), .Y(n8164) );
  OAI22X1 U6258 ( .A0(n3287), .A1(M2_mult_x_15_n43), .B0(n3288), .B1(n10388), 
        .Y(n10405) );
  NAND2BX1 U6259 ( .AN(n9700), .B(n3297), .Y(n3293) );
  INVXL U6260 ( .A(n12675), .Y(n3979) );
  INVX1 U6261 ( .A(n16151), .Y(n4128) );
  INVX1 U6262 ( .A(n16019), .Y(n3343) );
  NAND2X1 U6263 ( .A(n3744), .B(n12447), .Y(n3743) );
  OAI21XL U6264 ( .A0(n12706), .A1(n12707), .B0(n12705), .Y(n5998) );
  INVXL U6265 ( .A(n12706), .Y(n5999) );
  INVX1 U6266 ( .A(n12986), .Y(n12987) );
  NAND2X1 U6267 ( .A(n12790), .B(n12789), .Y(n12815) );
  NAND2BXL U6268 ( .AN(n9377), .B(n3269), .Y(n3267) );
  INVXL U6269 ( .A(n12380), .Y(n6136) );
  NAND2BXL U6270 ( .AN(n12134), .B(n3388), .Y(n3386) );
  OAI21XL U6271 ( .A0(n3287), .A1(n9617), .B0(n3302), .Y(n9618) );
  NAND2X1 U6272 ( .A(n4091), .B(n4193), .Y(n18359) );
  ADDFHX1 U6273 ( .A(n17612), .B(n17611), .CI(n17610), .CO(n17844), .S(n17643)
         );
  OAI2BB1XL U6274 ( .A0N(n17533), .A1N(n5862), .B0(n5861), .Y(n17577) );
  ADDFHX1 U6275 ( .A(n18459), .B(n18458), .CI(n18457), .CO(n18473), .S(n18514)
         );
  ADDFHX1 U6276 ( .A(n12158), .B(n12157), .CI(n12156), .CO(n12136), .S(n12214)
         );
  OAI22X1 U6277 ( .A0(n3287), .A1(n10169), .B0(n3288), .B1(n10309), .Y(n10315)
         );
  NAND2X1 U6278 ( .A(n17135), .B(n17134), .Y(n17378) );
  OR2XL U6279 ( .A(n10695), .B(n9161), .Y(n9160) );
  OAI2BB1XL U6280 ( .A0N(n17729), .A1N(n5795), .B0(n5793), .Y(n17759) );
  NAND2XL U6281 ( .A(n7179), .B(n7178), .Y(n3543) );
  NAND2XL U6282 ( .A(n12177), .B(n12176), .Y(n6003) );
  INVX1 U6283 ( .A(n7577), .Y(n5595) );
  OR2X2 U6284 ( .A(n9616), .B(n3288), .Y(n3302) );
  INVX1 U6285 ( .A(n11790), .Y(n4514) );
  OR2X2 U6286 ( .A(n12317), .B(n12316), .Y(n12260) );
  XNOR3X2 U6287 ( .A(n12104), .B(n3939), .C(n12103), .Y(n3388) );
  OAI21XL U6288 ( .A0(n4333), .A1(n3182), .B0(n4332), .Y(n9357) );
  ADDFHX1 U6289 ( .A(n12124), .B(n12123), .CI(n12122), .CO(n12134), .S(n12157)
         );
  NAND2X1 U6290 ( .A(n9159), .B(n10674), .Y(n9163) );
  XOR2X1 U6291 ( .A(n12177), .B(n12176), .Y(n4005) );
  AND2X2 U6292 ( .A(n21498), .B(n23398), .Y(n6189) );
  OR2X2 U6293 ( .A(n9402), .B(n3288), .Y(n3303) );
  ADDFHX2 U6294 ( .A(n18367), .B(n18366), .CI(n18365), .CO(n18360), .S(n18381)
         );
  XOR2X1 U6295 ( .A(n18549), .B(n5443), .Y(n18564) );
  INVXL U6296 ( .A(n6082), .Y(n6080) );
  NAND2X1 U6297 ( .A(n12805), .B(n12804), .Y(n12986) );
  AND2X1 U6298 ( .A(n18997), .B(n18996), .Y(n4704) );
  NAND2XL U6299 ( .A(n3498), .B(n3497), .Y(n6807) );
  NAND2X1 U6300 ( .A(n5564), .B(n5563), .Y(n7172) );
  INVX1 U6301 ( .A(n18996), .Y(n18714) );
  ADDFHX1 U6302 ( .A(n6886), .B(n6885), .CI(n6884), .CO(n6934), .S(n6897) );
  NAND2X1 U6303 ( .A(n14348), .B(n14347), .Y(n14678) );
  ADDFHX2 U6304 ( .A(n6386), .B(n6385), .CI(n6384), .CO(n6814), .S(n6387) );
  INVX8 U6305 ( .A(n3017), .Y(n3040) );
  OR2X2 U6306 ( .A(n10333), .B(n10403), .Y(n3290) );
  ADDFHX1 U6307 ( .A(n6996), .B(n6995), .CI(n6994), .CO(n7124), .S(n6998) );
  OR2XL U6308 ( .A(n11717), .B(n11716), .Y(n3645) );
  NAND2XL U6309 ( .A(n16120), .B(n16119), .Y(n3815) );
  OR2XL U6310 ( .A(n12311), .B(n12310), .Y(n12309) );
  NAND2XL U6311 ( .A(n16149), .B(n16148), .Y(n4831) );
  XOR2X1 U6312 ( .A(n16149), .B(n16148), .Y(n3847) );
  NAND2XL U6313 ( .A(n5777), .B(n3417), .Y(n5776) );
  OAI2BB1XL U6314 ( .A0N(n13791), .A1N(n13790), .B0(n25860), .Y(n13850) );
  NAND2X1 U6315 ( .A(n5424), .B(n5423), .Y(n18272) );
  ADDFHX2 U6316 ( .A(n16215), .B(n16214), .CI(n16213), .CO(n16259), .S(n16191)
         );
  INVX1 U6317 ( .A(n23124), .Y(n21444) );
  OAI21XL U6318 ( .A0(n16160), .A1(n16159), .B0(n16158), .Y(n5955) );
  NAND2BXL U6319 ( .AN(n11854), .B(n3915), .Y(n3914) );
  OR2X2 U6320 ( .A(n9317), .B(n10403), .Y(n3292) );
  NAND2XL U6321 ( .A(n12446), .B(n12445), .Y(n3745) );
  XOR2X1 U6322 ( .A(n11853), .B(n3916), .Y(n12434) );
  OAI2BB1X1 U6323 ( .A0N(n5669), .A1N(n16971), .B0(n5668), .Y(n16996) );
  NAND2X1 U6324 ( .A(n3041), .B(n19334), .Y(n19335) );
  NAND2XL U6325 ( .A(n3179), .B(n3953), .Y(n5691) );
  BUFX2 U6326 ( .A(n6778), .Y(n4769) );
  OR2X2 U6327 ( .A(n17151), .B(n17150), .Y(n17153) );
  OR2X2 U6328 ( .A(n12998), .B(n12997), .Y(n13000) );
  INVX1 U6329 ( .A(n6401), .Y(n3595) );
  OR2X2 U6330 ( .A(n14360), .B(n14359), .Y(n14362) );
  INVXL U6331 ( .A(n6400), .Y(n3517) );
  XOR2X1 U6332 ( .A(n18760), .B(n19029), .Y(n18769) );
  NAND2BXL U6333 ( .AN(n16091), .B(n3695), .Y(n3694) );
  AND2XL U6334 ( .A(n11854), .B(n3917), .Y(n3913) );
  XNOR2XL U6335 ( .A(n4808), .B(M2_mult_x_15_n1668), .Y(n10404) );
  INVX1 U6336 ( .A(n4745), .Y(n4746) );
  OR2XL U6337 ( .A(n18195), .B(n18194), .Y(n18193) );
  XNOR2X1 U6338 ( .A(n4565), .B(n3019), .Y(n4934) );
  OAI22X1 U6339 ( .A0(n3178), .A1(n9874), .B0(n10660), .B1(n9901), .Y(n4335)
         );
  INVX1 U6340 ( .A(n5980), .Y(n5982) );
  NAND2X1 U6341 ( .A(n23116), .B(n21405), .Y(n21396) );
  INVXL U6342 ( .A(n4739), .Y(n4740) );
  NAND2BX1 U6343 ( .AN(n4157), .B(n4156), .Y(n16000) );
  OAI21XL U6344 ( .A0(n12618), .A1(n3883), .B0(n4996), .Y(n11913) );
  OAI21X2 U6345 ( .A0(n8160), .A1(n8159), .B0(n8158), .Y(n8161) );
  NAND4X1 U6346 ( .A(n9124), .B(n9123), .C(n9122), .D(n25216), .Y(n10674) );
  INVX1 U6347 ( .A(M2_mult_x_15_n1668), .Y(n3177) );
  OAI22X1 U6348 ( .A0(n17964), .A1(n3195), .B0(n18483), .B1(n18467), .Y(n3440)
         );
  NAND2BXL U6349 ( .AN(n6975), .B(n3564), .Y(n3562) );
  INVXL U6350 ( .A(n3417), .Y(n3416) );
  NAND2XL U6351 ( .A(n16091), .B(n3697), .Y(n3693) );
  INVX8 U6352 ( .A(n19297), .Y(n3041) );
  BUFX8 U6353 ( .A(n12576), .Y(n12759) );
  NAND2BXL U6354 ( .AN(n7066), .B(n3541), .Y(n3540) );
  OAI22X1 U6355 ( .A0(n16977), .A1(n16048), .B0(n3105), .B1(n16047), .Y(n16091) );
  OAI22XL U6356 ( .A0(n12152), .A1(n12220), .B0(n3185), .B1(n6137), .Y(n12344)
         );
  INVXL U6357 ( .A(n3406), .Y(n3404) );
  OAI21XL U6358 ( .A0(n12598), .A1(n6008), .B0(n6007), .Y(n12155) );
  OAI22X1 U6359 ( .A0(n12597), .A1(n12165), .B0(n12595), .B1(n12126), .Y(
        n12154) );
  OAI21X2 U6360 ( .A0(n19289), .A1(n19288), .B0(n19287), .Y(n19290) );
  NAND4X1 U6361 ( .A(n14456), .B(n14444), .C(n14443), .D(n14442), .Y(n14712)
         );
  OAI22X1 U6362 ( .A0(n12003), .A1(n12715), .B0(n12525), .B1(n12002), .Y(n3417) );
  OAI22XL U6363 ( .A0(n16701), .A1(n6145), .B0(n16699), .B1(n16533), .Y(n16543) );
  OAI22X1 U6364 ( .A0(n3102), .A1(n16165), .B0(n16332), .B1(n16219), .Y(n16208) );
  NAND2X1 U6365 ( .A(n2978), .B(n4227), .Y(n4488) );
  NAND2BXL U6366 ( .AN(n7632), .B(n5122), .Y(n5109) );
  OAI22X1 U6367 ( .A0(n18242), .A1(n18052), .B0(n18168), .B1(n18027), .Y(
        n18064) );
  NOR2BXL U6368 ( .AN(n3110), .B(n16939), .Y(n16695) );
  XOR2X1 U6369 ( .A(n25884), .B(n3876), .Y(n3875) );
  AND2X2 U6370 ( .A(n12535), .B(n12995), .Y(n12996) );
  NAND2XL U6371 ( .A(n5770), .B(n20696), .Y(n4839) );
  NAND2XL U6372 ( .A(n21053), .B(n5770), .Y(n4838) );
  XOR2X1 U6373 ( .A(n25870), .B(n7800), .Y(n3451) );
  NAND2XL U6374 ( .A(n3792), .B(n3109), .Y(n3791) );
  OAI22X1 U6375 ( .A0(n17148), .A1(n3201), .B0(n3194), .B1(n3196), .Y(n17057)
         );
  CLKINVX3 U6376 ( .A(n5124), .Y(n3188) );
  OAI22X1 U6377 ( .A0(n3194), .A1(n3201), .B0(n17148), .B1(n3021), .Y(n17046)
         );
  XOR2X1 U6378 ( .A(M3_mult_x_15_b_1_), .B(n3755), .Y(n3754) );
  NAND2XL U6379 ( .A(n5770), .B(n21050), .Y(n4853) );
  NAND2XL U6380 ( .A(n20934), .B(n5770), .Y(n4854) );
  NAND2XL U6381 ( .A(n3790), .B(n3792), .Y(n3789) );
  NAND2X2 U6382 ( .A(n11749), .B(n5984), .Y(n12576) );
  NAND2XL U6383 ( .A(n4188), .B(M4_a_0_), .Y(n4187) );
  INVXL U6384 ( .A(n4592), .Y(n3541) );
  NOR2XL U6385 ( .A(n11728), .B(n12760), .Y(n3655) );
  OAI22XL U6386 ( .A0(n6323), .A1(n7288), .B0(n7287), .B1(n6364), .Y(n6383) );
  INVX8 U6387 ( .A(n3637), .Y(n16960) );
  XNOR2X1 U6388 ( .A(n3196), .B(n3022), .Y(n16922) );
  NAND2BXL U6389 ( .AN(n15965), .B(n3637), .Y(n3636) );
  OAI22X1 U6390 ( .A0(n17148), .A1(n3198), .B0(n3194), .B1(n3021), .Y(n16925)
         );
  AOI22XL U6391 ( .A0(n4566), .A1(data[18]), .B0(in_valid_d), .B1(w1[274]), 
        .Y(n9067) );
  AOI22XL U6392 ( .A0(n4566), .A1(data[16]), .B0(in_valid_d), .B1(w1[272]), 
        .Y(n9089) );
  BUFX3 U6393 ( .A(M1_a_9_), .Y(n4567) );
  NAND2X1 U6394 ( .A(n7978), .B(n8011), .Y(n8002) );
  AOI21X1 U6395 ( .A0(n8151), .A1(n8150), .B0(n8149), .Y(n8152) );
  INVX1 U6396 ( .A(n18226), .Y(n3192) );
  XOR2X1 U6397 ( .A(n12701), .B(n3903), .Y(n11642) );
  INVXL U6398 ( .A(n3413), .Y(n3371) );
  NAND2XL U6399 ( .A(n11658), .B(n5029), .Y(n5028) );
  NAND2BX1 U6400 ( .AN(n18223), .B(M4_U3_U1_or2_inv_0__30_), .Y(n3392) );
  BUFX3 U6401 ( .A(n12616), .Y(n12119) );
  XOR2X1 U6402 ( .A(n12225), .B(M3_mult_x_15_n1682), .Y(n12065) );
  AOI21XL U6403 ( .A0(n19145), .A1(n19144), .B0(n19143), .Y(n19146) );
  BUFX3 U6404 ( .A(M3_U3_U1_or2_inv_0__18_), .Y(n3903) );
  AND2X2 U6405 ( .A(n3111), .B(data[92]), .Y(n18754) );
  NOR2BXL U6406 ( .AN(n6944), .B(n7695), .Y(n6333) );
  NOR2X1 U6407 ( .A(n7989), .B(n8014), .Y(n8001) );
  XOR2X1 U6408 ( .A(n3201), .B(n6014), .Y(n16903) );
  AOI21X1 U6409 ( .A0(n14898), .A1(n14859), .B0(n14897), .Y(n14899) );
  NOR2XL U6410 ( .A(M4_a_2_), .B(n3206), .Y(M4_U3_U1_enc_tree_1__1__28_) );
  INVXL U6411 ( .A(M0_b_2_), .Y(n7057) );
  AND2XL U6412 ( .A(M0_U4_U1_or2_inv_0__18_), .B(n7621), .Y(n3529) );
  INVXL U6413 ( .A(n3376), .Y(M4_a_2_) );
  NOR2X1 U6414 ( .A(n8803), .B(n8298), .Y(n8125) );
  NAND2X1 U6415 ( .A(n3111), .B(sigma10[30]), .Y(n11551) );
  NOR2X1 U6416 ( .A(n8772), .B(n8308), .Y(n8116) );
  INVX1 U6417 ( .A(M5_a_22_), .Y(n15969) );
  BUFX12 U6418 ( .A(M3_mult_x_15_b_7_), .Y(n3197) );
  INVX1 U6419 ( .A(n16475), .Y(n3109) );
  OAI21XL U6420 ( .A0(n21288), .A1(n21287), .B0(n21286), .Y(n21289) );
  AOI21X1 U6421 ( .A0(n3223), .A1(sigma10[27]), .B0(n14412), .Y(n14705) );
  NOR2X1 U6422 ( .A(n8165), .B(n8184), .Y(n8110) );
  INVX1 U6423 ( .A(n3757), .Y(n3756) );
  OAI21XL U6424 ( .A0(n21234), .A1(n21233), .B0(n21232), .Y(n21291) );
  INVX1 U6425 ( .A(n25873), .Y(n7738) );
  AOI21XL U6426 ( .A0(n14789), .A1(n14788), .B0(n14787), .Y(n14790) );
  INVX4 U6427 ( .A(n25750), .Y(n3045) );
  NOR2X1 U6428 ( .A(n8067), .B(n8195), .Y(n8128) );
  INVX8 U6429 ( .A(n6326), .Y(n3046) );
  NOR2XL U6430 ( .A(n11294), .B(n11437), .Y(n11414) );
  NAND2XL U6431 ( .A(n25743), .B(y20[20]), .Y(n3601) );
  NOR2X1 U6432 ( .A(n8171), .B(n8203), .Y(n8138) );
  NOR2X1 U6433 ( .A(n8135), .B(n8199), .Y(n8086) );
  CLKINVX3 U6434 ( .A(n4789), .Y(n3213) );
  CLKINVX3 U6435 ( .A(M0_a_18_), .Y(n6281) );
  CLKINVX2 U6436 ( .A(n3216), .Y(n4573) );
  NOR2X1 U6437 ( .A(n19794), .B(n19392), .Y(n19178) );
  NOR2XL U6438 ( .A(n19551), .B(n19537), .Y(n19139) );
  OAI2BB1X1 U6439 ( .A0N(y10[26]), .A1N(n3224), .B0(n7396), .Y(n7857) );
  CLKINVX2 U6440 ( .A(n3216), .Y(n4574) );
  CLKINVX2 U6441 ( .A(n3216), .Y(n4572) );
  NOR2XL U6442 ( .A(n19479), .B(n19385), .Y(n19175) );
  CLKINVX2 U6443 ( .A(n3216), .Y(n4571) );
  BUFX3 U6444 ( .A(n25741), .Y(n20890) );
  NAND2X1 U6445 ( .A(n4856), .B(target_temp[30]), .Y(n14405) );
  OAI2BB1XL U6446 ( .A0N(y12[30]), .A1N(n4856), .B0(n9110), .Y(n9113) );
  INVX8 U6447 ( .A(n16631), .Y(n3047) );
  NOR2X1 U6448 ( .A(n19212), .B(n19254), .Y(n19219) );
  NAND3X1 U6449 ( .A(n11587), .B(n11586), .C(n11585), .Y(n18786) );
  OAI2BB1X2 U6450 ( .A0N(n3758), .A1N(data[80]), .B0(n17475), .Y(n3757) );
  AND2X2 U6451 ( .A(n5016), .B(n5013), .Y(n4663) );
  XNOR2X1 U6452 ( .A(n7621), .B(n25869), .Y(n3542) );
  NOR2X1 U6453 ( .A(n19815), .B(n19370), .Y(n19170) );
  AOI222XL U6454 ( .A0(n22928), .A1(n26493), .B0(n22700), .B1(n11059), .C0(
        n22927), .C1(n11058), .Y(n22929) );
  NOR2BX2 U6455 ( .AN(n4101), .B(n2987), .Y(n5729) );
  CLKINVX3 U6456 ( .A(M0_a_3_), .Y(n6989) );
  NAND3X1 U6457 ( .A(n11595), .B(n11594), .C(n11593), .Y(n18776) );
  INVX1 U6458 ( .A(n8355), .Y(n8378) );
  CLKBUFX2 U6459 ( .A(n22897), .Y(n10797) );
  NOR2X1 U6460 ( .A(n15942), .B(n25912), .Y(n4539) );
  NOR2X1 U6461 ( .A(n14917), .B(n14950), .Y(n14887) );
  AOI22X1 U6462 ( .A0(n5770), .A1(data[72]), .B0(w2[40]), .B1(in_valid_t), .Y(
        n4520) );
  NAND4X1 U6463 ( .A(n7964), .B(n7963), .C(n7962), .D(n7961), .Y(n8256) );
  CLKINVX3 U6464 ( .A(n3117), .Y(n3113) );
  NAND2XL U6465 ( .A(n5480), .B(sigma11[5]), .Y(n5891) );
  OAI22X1 U6466 ( .A0(n15941), .A1(n6186), .B0(n15940), .B1(n23988), .Y(n4536)
         );
  NAND4X1 U6467 ( .A(n7940), .B(n7939), .C(n7938), .D(n7937), .Y(n8357) );
  NAND2XL U6468 ( .A(n5480), .B(sigma11[12]), .Y(n5872) );
  INVXL U6469 ( .A(n25796), .Y(n3758) );
  NAND4X1 U6470 ( .A(n7982), .B(n7981), .C(n7980), .D(n7979), .Y(n8235) );
  OAI22XL U6471 ( .A0(n15942), .A1(n26516), .B0(n26033), .B1(n17167), .Y(n4534) );
  NAND4X1 U6472 ( .A(n7975), .B(n7974), .C(n7973), .D(n7972), .Y(n8261) );
  OAI22X4 U6473 ( .A0(n6207), .A1(n4860), .B0(n25911), .B1(n25796), .Y(n11495)
         );
  NOR2X1 U6474 ( .A(n15557), .B(n15052), .Y(n14838) );
  OR2XL U6475 ( .A(n3115), .B(n23980), .Y(n9153) );
  BUFX8 U6476 ( .A(n25229), .Y(n4856) );
  NOR2X1 U6477 ( .A(n15413), .B(n15005), .Y(n14798) );
  NOR2X1 U6478 ( .A(n15422), .B(n14980), .Y(n14745) );
  CLKINVX4 U6479 ( .A(n26491), .Y(n3217) );
  CLKINVX4 U6480 ( .A(n22549), .Y(n23109) );
  NOR2XL U6481 ( .A(n21228), .B(n21212), .Y(n21231) );
  CLKINVX4 U6482 ( .A(n26490), .Y(n3219) );
  AND2X2 U6483 ( .A(n6232), .B(n3585), .Y(n3584) );
  OAI22X1 U6484 ( .A0(n25796), .A1(n26262), .B0(n26015), .B1(n15940), .Y(n4921) );
  NOR2X1 U6485 ( .A(n15547), .B(n15047), .Y(n14832) );
  NAND2X1 U6486 ( .A(n25229), .B(target_temp[17]), .Y(n13356) );
  NOR2X1 U6487 ( .A(n21325), .B(n21370), .Y(n21326) );
  NOR2X1 U6488 ( .A(n25796), .B(n25886), .Y(n25201) );
  NAND2X1 U6489 ( .A(n25229), .B(target_temp[18]), .Y(n11537) );
  INVX1 U6490 ( .A(n19390), .Y(n19787) );
  NAND2XL U6491 ( .A(n25229), .B(y12[14]), .Y(n5762) );
  NOR2X1 U6492 ( .A(n21301), .B(n21341), .Y(n21302) );
  NOR2X1 U6493 ( .A(n15435), .B(n14986), .Y(n14749) );
  NOR2X1 U6494 ( .A(n15461), .B(n15056), .Y(n14821) );
  AOI22X1 U6495 ( .A0(n5480), .A1(sigma11[20]), .B0(in_valid_t), .B1(w2[52]), 
        .Y(n17477) );
  NAND2X1 U6496 ( .A(n3120), .B(y20[27]), .Y(n8087) );
  NOR2XL U6497 ( .A(n21201), .B(n21626), .Y(n21204) );
  NAND2X1 U6498 ( .A(n3120), .B(y20[28]), .Y(n8099) );
  NOR2XL U6499 ( .A(n21220), .B(n21554), .Y(n21223) );
  INVX1 U6500 ( .A(n15103), .Y(n15126) );
  XNOR2X1 U6501 ( .A(n3119), .B(n11210), .Y(n21057) );
  BUFX3 U6502 ( .A(n23089), .Y(n9109) );
  INVX1 U6503 ( .A(n14996), .Y(n15075) );
  NOR2XL U6504 ( .A(n21261), .B(n21473), .Y(n21264) );
  NAND2X1 U6505 ( .A(n3120), .B(y20[23]), .Y(n8061) );
  CLKINVX3 U6506 ( .A(n3225), .Y(n3116) );
  BUFX2 U6507 ( .A(n11146), .Y(n11073) );
  NAND2X1 U6508 ( .A(n3120), .B(y20[26]), .Y(n8092) );
  BUFX2 U6509 ( .A(n11144), .Y(n11063) );
  CLKINVX8 U6510 ( .A(n3024), .Y(n3050) );
  AOI21XL U6511 ( .A0(n4718), .A1(n21166), .B0(n4980), .Y(n4969) );
  AOI21X1 U6512 ( .A0(n21166), .A1(n4717), .B0(n5987), .Y(n5986) );
  INVX1 U6513 ( .A(n15155), .Y(n15169) );
  NOR2XL U6514 ( .A(n21225), .B(n21469), .Y(n21228) );
  XOR2X2 U6515 ( .A(n23170), .B(n23169), .Y(n23955) );
  AND2X2 U6516 ( .A(n21379), .B(n21413), .Y(n21382) );
  INVX8 U6517 ( .A(n11479), .Y(n25796) );
  NOR2XL U6518 ( .A(n21371), .B(n21405), .Y(n21320) );
  INVX4 U6519 ( .A(n23039), .Y(n23428) );
  INVX4 U6520 ( .A(n23133), .Y(n23429) );
  INVX8 U6521 ( .A(n3226), .Y(n25541) );
  INVXL U6522 ( .A(n21616), .Y(n21219) );
  BUFX2 U6523 ( .A(n11154), .Y(n11059) );
  BUFX2 U6524 ( .A(n11152), .Y(n11058) );
  OAI21X1 U6525 ( .A0(n14833), .A1(n26514), .B0(n8103), .Y(n8184) );
  OAI21X1 U6526 ( .A0(n14833), .A1(n23789), .B0(n8085), .Y(n8203) );
  OAI21XL U6527 ( .A0(n14833), .A1(n26190), .B0(n14846), .Y(n14927) );
  BUFX2 U6528 ( .A(n11163), .Y(n10749) );
  OAI21X1 U6529 ( .A0(n14833), .A1(n26545), .B0(n8080), .Y(n8199) );
  CLKINVX2 U6530 ( .A(n11168), .Y(n3225) );
  OAI21X1 U6531 ( .A0(n19237), .A1(n14966), .B0(n14965), .Y(n23169) );
  OAI22X1 U6532 ( .A0(n23193), .A1(n26231), .B0(n9107), .B1(n25938), .Y(n11140) );
  CLKINVX3 U6533 ( .A(n26489), .Y(n3119) );
  NOR2X1 U6534 ( .A(n7382), .B(n26045), .Y(n7378) );
  INVXL U6535 ( .A(n11220), .Y(n22621) );
  AOI22X1 U6536 ( .A0(n3027), .A1(w2[57]), .B0(n19216), .B1(w1[89]), .Y(n19223) );
  INVX8 U6537 ( .A(n25696), .Y(n3057) );
  AND2X1 U6538 ( .A(n2982), .B(temp2[30]), .Y(n4712) );
  AOI22XL U6539 ( .A0(n19216), .A1(w1[110]), .B0(n19346), .B1(w2[78]), .Y(
        n4466) );
  INVX2 U6540 ( .A(n25856), .Y(n23985) );
  AOI22X1 U6541 ( .A0(w2[87]), .A1(n19349), .B0(n3026), .B1(w1[119]), .Y(
        n14834) );
  NAND2X1 U6542 ( .A(n3027), .B(w2[23]), .Y(n8063) );
  XNOR2X1 U6543 ( .A(n11210), .B(n11169), .Y(n11090) );
  OR2XL U6544 ( .A(n21195), .B(n21623), .Y(n21189) );
  AOI22X1 U6545 ( .A0(y10[29]), .A1(n19235), .B0(n3026), .B1(temp1[29]), .Y(
        n8109) );
  INVX4 U6546 ( .A(n25693), .Y(n3060) );
  INVX1 U6547 ( .A(n25664), .Y(n3227) );
  BUFX3 U6548 ( .A(n9108), .Y(n11311) );
  NAND2X1 U6549 ( .A(n11194), .B(n11193), .Y(n21089) );
  INVX8 U6550 ( .A(n4637), .Y(n19237) );
  NAND2X1 U6551 ( .A(n11088), .B(n11087), .Y(n11169) );
  INVX4 U6552 ( .A(n21111), .Y(n3062) );
  INVX8 U6553 ( .A(n4637), .Y(n3063) );
  NOR2X1 U6554 ( .A(n17167), .B(n24000), .Y(n6155) );
  INVX1 U6555 ( .A(valid[0]), .Y(n3501) );
  INVX1 U6556 ( .A(n25143), .Y(n9062) );
  INVX1 U6557 ( .A(n25153), .Y(n9045) );
  INVX2 U6558 ( .A(n25149), .Y(n5567) );
  NAND2X1 U6559 ( .A(in_valid_t), .B(learning_rate[28]), .Y(n11581) );
  NOR2XL U6560 ( .A(n15940), .B(n26005), .Y(n4980) );
  NAND2X1 U6561 ( .A(in_valid_t), .B(w2[41]), .Y(n4661) );
  NAND2X1 U6562 ( .A(in_valid_t), .B(w2[42]), .Y(n4660) );
  AND2X2 U6563 ( .A(in_valid_t), .B(w2[47]), .Y(n4654) );
  NOR2XL U6564 ( .A(n15940), .B(n26016), .Y(n4538) );
  NOR2XL U6565 ( .A(n15940), .B(n26006), .Y(n4896) );
  NOR2XL U6566 ( .A(n15940), .B(n26040), .Y(n4530) );
  NOR2X1 U6567 ( .A(n15940), .B(n26014), .Y(n5420) );
  NOR2XL U6568 ( .A(n15940), .B(n25997), .Y(n3982) );
  INVX8 U6569 ( .A(n4581), .Y(n4579) );
  NOR2X1 U6570 ( .A(n4583), .B(in_valid_w1), .Y(n25848) );
  INVX1 U6571 ( .A(data_point[3]), .Y(n6235) );
  INVX1 U6572 ( .A(data_point[4]), .Y(n6260) );
  INVX1 U6573 ( .A(data_point[6]), .Y(n6244) );
  INVX1 U6574 ( .A(data_point[0]), .Y(n6229) );
  INVXL U6575 ( .A(n4582), .Y(n3066) );
  AOI21XL U6576 ( .A0(n19089), .A1(n24525), .B0(n24486), .Y(n2397) );
  AOI22XL U6577 ( .A0(n24692), .A1(n25003), .B0(n24908), .B1(n25002), .Y(
        n25004) );
  INVX1 U6578 ( .A(n24631), .Y(n25508) );
  AOI21X1 U6579 ( .A0(n3602), .A1(n25744), .B0(n3600), .Y(n2380) );
  XOR2X1 U6580 ( .A(n24763), .B(n24762), .Y(n24764) );
  INVX1 U6581 ( .A(n24479), .Y(n25609) );
  AOI22X1 U6582 ( .A0(n3029), .A1(n24663), .B0(n25290), .B1(n24662), .Y(n25497) );
  AOI22X1 U6583 ( .A0(n3029), .A1(n24507), .B0(n25290), .B1(n24506), .Y(n25598) );
  AOI22X1 U6584 ( .A0(n3029), .A1(n24637), .B0(n25290), .B1(n24636), .Y(n25510) );
  INVX1 U6585 ( .A(n20684), .Y(n25623) );
  AOI22X1 U6586 ( .A0(n3029), .A1(n24670), .B0(n25290), .B1(n24669), .Y(n25487) );
  AOI22X1 U6587 ( .A0(n3029), .A1(n24518), .B0(n25290), .B1(n24517), .Y(n25579) );
  AOI22X1 U6588 ( .A0(n3029), .A1(n24780), .B0(n25290), .B1(n24779), .Y(n25449) );
  AOI22X1 U6589 ( .A0(n3029), .A1(n24771), .B0(n25290), .B1(n15906), .Y(n25461) );
  AOI22X1 U6590 ( .A0(n3029), .A1(n24502), .B0(n25290), .B1(n24484), .Y(n25611) );
  INVX1 U6591 ( .A(n24598), .Y(n25533) );
  AOI22X1 U6592 ( .A0(n3029), .A1(n25024), .B0(n25290), .B1(n25023), .Y(n25373) );
  AOI22X1 U6593 ( .A0(n3029), .A1(n24880), .B0(n25290), .B1(n21014), .Y(n25423) );
  AOI22X1 U6594 ( .A0(n3029), .A1(n24618), .B0(n25290), .B1(n24603), .Y(n25536) );
  AOI22X1 U6595 ( .A0(n3029), .A1(n24541), .B0(n25290), .B1(n24540), .Y(n25569) );
  AOI22X1 U6596 ( .A0(n3029), .A1(n24974), .B0(n25290), .B1(n24932), .Y(n25394) );
  AOI22X1 U6597 ( .A0(n3029), .A1(n24980), .B0(n25290), .B1(n24979), .Y(n25386) );
  XOR2X1 U6598 ( .A(n24609), .B(n24608), .Y(n24610) );
  INVX1 U6599 ( .A(n25323), .Y(n25732) );
  XOR2X1 U6600 ( .A(n24649), .B(n24648), .Y(n24650) );
  XOR2X1 U6601 ( .A(n24628), .B(n24645), .Y(n24629) );
  AOI21XL U6602 ( .A0(n24548), .A1(n25675), .B0(n24547), .Y(n2402) );
  INVX1 U6603 ( .A(n23720), .Y(n25422) );
  XNOR2X1 U6604 ( .A(n25358), .B(n24815), .Y(n24816) );
  INVX1 U6605 ( .A(n23841), .Y(n25385) );
  AOI222XL U6606 ( .A0(n23758), .A1(n25737), .B0(n25743), .B1(y20[16]), .C0(
        n25436), .C1(n20890), .Y(n2376) );
  INVX1 U6607 ( .A(n25826), .Y(n25824) );
  AOI21X1 U6608 ( .A0(n24743), .A1(n3060), .B0(n24742), .Y(n2420) );
  INVX1 U6609 ( .A(n23756), .Y(n25436) );
  OAI21XL U6610 ( .A0(n24419), .A1(n3057), .B0(n24418), .Y(n24420) );
  OAI21XL U6611 ( .A0(n23695), .A1(n3057), .B0(n23694), .Y(n23696) );
  INVX1 U6612 ( .A(n24488), .Y(n25610) );
  INVX1 U6613 ( .A(n24546), .Y(n25568) );
  INVX1 U6614 ( .A(n25689), .Y(n25742) );
  INVX1 U6615 ( .A(n23699), .Y(n25546) );
  XOR2X1 U6616 ( .A(n21013), .B(n21012), .Y(n21014) );
  INVX1 U6617 ( .A(n24473), .Y(n25624) );
  OAI21XL U6618 ( .A0(n24423), .A1(n3227), .B0(n24422), .Y(n24424) );
  INVX1 U6619 ( .A(n23768), .Y(n25535) );
  INVX1 U6620 ( .A(n25308), .Y(n25739) );
  INVX1 U6621 ( .A(n24523), .Y(n25578) );
  INVX1 U6622 ( .A(n24512), .Y(n25597) );
  XOR2X1 U6623 ( .A(n24701), .B(n24700), .Y(n24702) );
  OAI21XL U6624 ( .A0(n23877), .A1(n3227), .B0(n23876), .Y(n23878) );
  NAND2X1 U6625 ( .A(n24812), .B(n24811), .Y(n24814) );
  INVX1 U6626 ( .A(n24317), .Y(n24325) );
  AOI22X1 U6627 ( .A0(n20385), .A1(n20918), .B0(n25300), .B1(n20917), .Y(
        n24488) );
  XNOR2X1 U6628 ( .A(n24550), .B(n24549), .Y(n24551) );
  XNOR2X1 U6629 ( .A(n24529), .B(n24528), .Y(n24530) );
  INVX1 U6630 ( .A(n25103), .Y(n25113) );
  XOR2X1 U6631 ( .A(n23831), .B(n23830), .Y(n23832) );
  AOI22X1 U6632 ( .A0(n20385), .A1(n23625), .B0(n25300), .B1(n23624), .Y(
        n24546) );
  XOR2X1 U6633 ( .A(n23803), .B(n23802), .Y(n23804) );
  INVX1 U6634 ( .A(n24405), .Y(n24456) );
  AOI22X1 U6635 ( .A0(n20385), .A1(n20898), .B0(n25300), .B1(n20897), .Y(
        n24523) );
  INVX1 U6636 ( .A(n25853), .Y(n25845) );
  XOR2X1 U6637 ( .A(n24620), .B(n24619), .Y(n24621) );
  INVX1 U6638 ( .A(n25095), .Y(n25083) );
  AOI22X1 U6639 ( .A0(n20385), .A1(n24566), .B0(n25300), .B1(n24565), .Y(
        n25308) );
  XOR2X1 U6640 ( .A(n24635), .B(n24657), .Y(n24636) );
  OAI21X1 U6641 ( .A0(n4788), .A1(n23813), .B0(n23812), .Y(n24421) );
  OAI21X1 U6642 ( .A0(n4788), .A1(n23819), .B0(n23818), .Y(n24417) );
  XNOR2X1 U6643 ( .A(n24539), .B(n24538), .Y(n24540) );
  XNOR2X1 U6644 ( .A(n24589), .B(n24588), .Y(n24590) );
  XOR2X1 U6645 ( .A(n24710), .B(n24709), .Y(n24711) );
  OAI21X1 U6646 ( .A0(n4788), .A1(n23693), .B0(n23692), .Y(n25801) );
  AOI222X1 U6647 ( .A0(n4791), .A1(n24430), .B0(n24292), .B1(n24428), .C0(
        n24427), .C1(n24291), .Y(n25095) );
  XNOR2X1 U6648 ( .A(n23829), .B(n23752), .Y(n23753) );
  INVX4 U6649 ( .A(n15818), .Y(n25290) );
  NAND2X1 U6650 ( .A(n24428), .B(n24059), .Y(n4450) );
  XOR2X1 U6651 ( .A(n20904), .B(n20903), .Y(n20905) );
  OAI21X1 U6652 ( .A0(n4788), .A1(n23875), .B0(n23874), .Y(n25712) );
  AOI222X1 U6653 ( .A0(n24431), .A1(n24430), .B0(n24429), .B1(n24428), .C0(
        n24427), .C1(n24426), .Y(n25103) );
  AOI222X1 U6654 ( .A0(n4793), .A1(n24430), .B0(n24400), .B1(n24428), .C0(
        n24427), .C1(n24399), .Y(n24405) );
  XOR2X1 U6655 ( .A(n20875), .B(n20874), .Y(n20876) );
  XNOR2X1 U6656 ( .A(n24493), .B(n24477), .Y(n24478) );
  NAND2X1 U6657 ( .A(n15934), .B(n24667), .Y(n15936) );
  XNOR2X1 U6658 ( .A(n20887), .B(n20886), .Y(n20888) );
  INVX1 U6659 ( .A(n20994), .Y(n24572) );
  AND4X4 U6660 ( .A(n20384), .B(n20383), .C(n20382), .D(n20425), .Y(n20385) );
  NOR2X2 U6661 ( .A(n24071), .B(n24070), .Y(n24434) );
  NOR2X1 U6662 ( .A(n24977), .B(n24976), .Y(n25284) );
  NOR2X1 U6663 ( .A(n24569), .B(n20227), .Y(n20234) );
  XOR2X1 U6664 ( .A(n24505), .B(n24504), .Y(n24506) );
  XNOR2X1 U6665 ( .A(n23623), .B(n23622), .Y(n23624) );
  AOI222XL U6666 ( .A0(n23249), .A1(n23429), .B0(n23428), .B1(target_temp[10]), 
        .C0(in_valid_t), .C1(target[10]), .Y(n2242) );
  AOI222XL U6667 ( .A0(n23353), .A1(n23429), .B0(n23428), .B1(target_temp[6]), 
        .C0(in_valid_t), .C1(target[6]), .Y(n2238) );
  AOI222XL U6668 ( .A0(n23357), .A1(n23429), .B0(n23428), .B1(target_temp[7]), 
        .C0(in_valid_t), .C1(target[7]), .Y(n2239) );
  AOI222XL U6669 ( .A0(n23354), .A1(n23429), .B0(n23428), .B1(target_temp[5]), 
        .C0(in_valid_t), .C1(target[5]), .Y(n2237) );
  AOI222XL U6670 ( .A0(n23352), .A1(n23429), .B0(n23428), .B1(target_temp[8]), 
        .C0(in_valid_t), .C1(target[8]), .Y(n2240) );
  AOI222XL U6671 ( .A0(n23361), .A1(n23429), .B0(n23428), .B1(target_temp[11]), 
        .C0(in_valid_t), .C1(target[11]), .Y(n2243) );
  AOI222XL U6672 ( .A0(n23390), .A1(n23429), .B0(n23428), .B1(target_temp[19]), 
        .C0(in_valid_t), .C1(target[19]), .Y(n2251) );
  AOI222XL U6673 ( .A0(n23358), .A1(n23429), .B0(n23428), .B1(target_temp[17]), 
        .C0(in_valid_t), .C1(target[17]), .Y(n2249) );
  AOI222XL U6674 ( .A0(n23248), .A1(n23429), .B0(n23428), .B1(target_temp[9]), 
        .C0(in_valid_t), .C1(target[9]), .Y(n2241) );
  AOI222XL U6675 ( .A0(n23360), .A1(n23429), .B0(n23428), .B1(target_temp[12]), 
        .C0(in_valid_t), .C1(target[12]), .Y(n2244) );
  AOI222XL U6676 ( .A0(n23364), .A1(n23429), .B0(n23428), .B1(target_temp[2]), 
        .C0(in_valid_t), .C1(target[2]), .Y(n2234) );
  AOI222XL U6677 ( .A0(n23365), .A1(n23429), .B0(n23428), .B1(target_temp[3]), 
        .C0(in_valid_t), .C1(target[3]), .Y(n2235) );
  AOI222XL U6678 ( .A0(n23362), .A1(n23429), .B0(n23428), .B1(target_temp[18]), 
        .C0(in_valid_t), .C1(target[18]), .Y(n2250) );
  AOI222XL U6679 ( .A0(n23359), .A1(n23429), .B0(n23428), .B1(target_temp[15]), 
        .C0(in_valid_t), .C1(target[15]), .Y(n2247) );
  AOI222XL U6680 ( .A0(n23368), .A1(n23429), .B0(n23428), .B1(target_temp[13]), 
        .C0(in_valid_t), .C1(target[13]), .Y(n2245) );
  AOI222XL U6681 ( .A0(n23367), .A1(n23429), .B0(n23428), .B1(target_temp[14]), 
        .C0(in_valid_t), .C1(target[14]), .Y(n2246) );
  AOI222XL U6682 ( .A0(n23363), .A1(n23429), .B0(n23428), .B1(target_temp[1]), 
        .C0(in_valid_t), .C1(target[1]), .Y(n2233) );
  AOI222XL U6683 ( .A0(n23389), .A1(n23429), .B0(n23428), .B1(target_temp[20]), 
        .C0(in_valid_t), .C1(target[20]), .Y(n2252) );
  AOI222XL U6684 ( .A0(n23391), .A1(n23429), .B0(n23428), .B1(target_temp[21]), 
        .C0(in_valid_t), .C1(target[21]), .Y(n2253) );
  AOI222XL U6685 ( .A0(n23366), .A1(n23429), .B0(n23428), .B1(target_temp[16]), 
        .C0(in_valid_t), .C1(target[16]), .Y(n2248) );
  AND3X2 U6686 ( .A(n20384), .B(n23175), .C(n9034), .Y(n4621) );
  NOR2X1 U6687 ( .A(n24583), .B(n15897), .Y(n15902) );
  AOI22XL U6688 ( .A0(n23256), .A1(n23387), .B0(n23257), .B1(n23386), .Y(
        n23388) );
  AOI22XL U6689 ( .A0(n23256), .A1(n23380), .B0(n23257), .B1(n23379), .Y(
        n23381) );
  AOI22XL U6690 ( .A0(n23256), .A1(n23376), .B0(n23257), .B1(n23327), .Y(
        n23328) );
  AOI22XL U6691 ( .A0(n23256), .A1(n23374), .B0(n23257), .B1(n23373), .Y(
        n23375) );
  NOR2X1 U6692 ( .A(n23827), .B(n20575), .Y(n23798) );
  AOI22XL U6693 ( .A0(n23256), .A1(n23305), .B0(n23257), .B1(n23304), .Y(
        n23306) );
  AOI22XL U6694 ( .A0(n23256), .A1(n23242), .B0(n23257), .B1(n23241), .Y(
        n23243) );
  AOI22XL U6695 ( .A0(n23256), .A1(n23290), .B0(n23257), .B1(n23289), .Y(
        n23291) );
  AOI22XL U6696 ( .A0(n23256), .A1(n23270), .B0(n23257), .B1(n23269), .Y(
        n23271) );
  AOI22XL U6697 ( .A0(n23256), .A1(n23275), .B0(n23257), .B1(n23274), .Y(
        n23276) );
  AOI22XL U6698 ( .A0(n23256), .A1(n23272), .B0(n23257), .B1(n23258), .Y(
        n23355) );
  AOI22XL U6699 ( .A0(n23256), .A1(n23277), .B0(n23257), .B1(n23252), .Y(
        n23324) );
  AOI22XL U6700 ( .A0(n23256), .A1(n23285), .B0(n23257), .B1(n23284), .Y(
        n23286) );
  AOI22XL U6701 ( .A0(n23256), .A1(n23297), .B0(n23257), .B1(n23296), .Y(
        n23298) );
  AOI22XL U6702 ( .A0(n23256), .A1(n23265), .B0(n23257), .B1(n23264), .Y(
        n23266) );
  AOI22XL U6703 ( .A0(n23256), .A1(n23318), .B0(n23257), .B1(n23246), .Y(
        n23247) );
  XOR2X1 U6704 ( .A(n20911), .B(n20910), .Y(n20912) );
  AOI22XL U6705 ( .A0(n23256), .A1(n23322), .B0(n23257), .B1(n23321), .Y(
        n23323) );
  AOI22XL U6706 ( .A0(n23256), .A1(n23316), .B0(n23257), .B1(n23315), .Y(
        n23317) );
  AOI22XL U6707 ( .A0(n23256), .A1(n23282), .B0(n23257), .B1(n23281), .Y(
        n23283) );
  AOI22XL U6708 ( .A0(n23256), .A1(n23350), .B0(n23257), .B1(n23349), .Y(
        n23351) );
  NOR2X1 U6709 ( .A(n24561), .B(n20523), .Y(n20528) );
  AOI22XL U6710 ( .A0(n23256), .A1(n23311), .B0(n23257), .B1(n23310), .Y(
        n23312) );
  AOI22XL U6711 ( .A0(n23256), .A1(n23335), .B0(n23257), .B1(n23334), .Y(
        n23336) );
  INVX1 U6712 ( .A(n24881), .Y(n4781) );
  AOI22XL U6713 ( .A0(n23256), .A1(n23341), .B0(n23257), .B1(n23340), .Y(
        n23342) );
  AOI222XL U6714 ( .A0(n23427), .A1(n3216), .B0(n4578), .B1(w1[280]), .C0(
        n25567), .C1(w1[312]), .Y(n2107) );
  AOI222XL U6715 ( .A0(n23426), .A1(n3216), .B0(n4577), .B1(w1[285]), .C0(
        n25567), .C1(w1[317]), .Y(n2127) );
  AOI222XL U6716 ( .A0(n23424), .A1(n3216), .B0(n21113), .B1(w1[284]), .C0(
        n25567), .C1(w1[316]), .Y(n2123) );
  AOI222XL U6717 ( .A0(n23422), .A1(n3216), .B0(n4576), .B1(w1[282]), .C0(
        n25567), .C1(w1[314]), .Y(n2115) );
  AOI222XL U6718 ( .A0(n23430), .A1(n3216), .B0(n4578), .B1(w1[281]), .C0(
        n25567), .C1(w1[313]), .Y(n2111) );
  INVX1 U6719 ( .A(n20635), .Y(n23799) );
  AOI222XL U6720 ( .A0(n23425), .A1(n3216), .B0(n4577), .B1(w1[279]), .C0(
        n23088), .C1(w1[311]), .Y(n2103) );
  INVX1 U6721 ( .A(n15751), .Y(n4452) );
  XOR2X1 U6722 ( .A(n23378), .B(n23377), .Y(n23379) );
  NAND2X1 U6723 ( .A(n4443), .B(n15748), .Y(n15750) );
  XOR2X1 U6724 ( .A(n23333), .B(n23332), .Y(n23334) );
  XOR2X1 U6725 ( .A(n23303), .B(n23302), .Y(n23304) );
  XOR2X1 U6726 ( .A(n23385), .B(n23384), .Y(n23386) );
  AOI21X1 U6727 ( .A0(n20556), .A1(n20576), .B0(n20509), .Y(n20906) );
  XOR2X1 U6728 ( .A(n23348), .B(n23347), .Y(n23349) );
  OAI22XL U6729 ( .A0(n15854), .A1(n3125), .B0(n15851), .B1(n15808), .Y(n15891) );
  XOR2X1 U6730 ( .A(n23320), .B(n23319), .Y(n23321) );
  AOI222X1 U6731 ( .A0(n23413), .A1(n23419), .B0(n23418), .B1(n23412), .C0(
        n23411), .C1(n23415), .Y(n23414) );
  XNOR2X1 U6732 ( .A(n23383), .B(n23326), .Y(n23327) );
  XNOR2X1 U6733 ( .A(n23263), .B(n23262), .Y(n23264) );
  XNOR2X1 U6734 ( .A(n23346), .B(n23245), .Y(n23246) );
  NAND2X1 U6735 ( .A(n20148), .B(n3032), .Y(n20228) );
  NAND3BX1 U6736 ( .AN(n15763), .B(n15815), .C(n15762), .Y(n15770) );
  XNOR2X1 U6737 ( .A(n23240), .B(n23239), .Y(n23241) );
  NAND2X1 U6738 ( .A(n15858), .B(n3125), .Y(n15894) );
  AOI2BB2X1 U6739 ( .B0(n23691), .B1(n8991), .A0N(n8991), .A1N(n23691), .Y(
        n23689) );
  NOR2X1 U6740 ( .A(n20179), .B(n20178), .Y(n20213) );
  INVX1 U6741 ( .A(n23237), .Y(n23293) );
  NAND2X1 U6742 ( .A(n3030), .B(n24063), .Y(n20152) );
  XNOR2X1 U6743 ( .A(n23278), .B(n23251), .Y(n23252) );
  AOI2BB2XL U6744 ( .B0(n8984), .B1(n8983), .A0N(n8983), .A1N(n8984), .Y(n9029) );
  NOR2BXL U6745 ( .AN(n20496), .B(n20473), .Y(n20526) );
  NOR2X1 U6746 ( .A(n15882), .B(n15808), .Y(n15849) );
  AND3X1 U6747 ( .A(n25274), .B(n25273), .C(n25272), .Y(n6219) );
  NOR2X1 U6748 ( .A(n15813), .B(n15812), .Y(n15846) );
  OAI21X2 U6749 ( .A0(n23224), .A1(n22215), .B0(n22214), .Y(n23228) );
  NOR2X1 U6750 ( .A(n23261), .B(n22391), .Y(n22408) );
  NOR2X1 U6751 ( .A(n25271), .B(n15705), .Y(n15766) );
  NAND2X1 U6752 ( .A(n23290), .B(n23287), .Y(n23250) );
  NAND2XL U6753 ( .A(n24309), .B(n20125), .Y(n20126) );
  NOR2X1 U6754 ( .A(n23267), .B(n23268), .Y(n23287) );
  NAND2BX2 U6755 ( .AN(n22184), .B(n6212), .Y(n23226) );
  OR3X2 U6756 ( .A(n23396), .B(n23411), .C(n22183), .Y(n6212) );
  INVX8 U6757 ( .A(n3124), .Y(n3067) );
  AND2X1 U6758 ( .A(n22389), .B(n22124), .Y(n6188) );
  NAND3BX1 U6759 ( .AN(n22195), .B(n22268), .C(n22194), .Y(n22200) );
  INVX1 U6760 ( .A(n22181), .Y(n23232) );
  OAI2BB1X2 U6761 ( .A0N(n15716), .A1N(n15717), .B0(n3133), .Y(n4456) );
  NOR3X1 U6762 ( .A(n23216), .B(n23215), .C(n23214), .Y(n25665) );
  AOI22X1 U6763 ( .A0(n22396), .A1(n3129), .B0(n22426), .B1(n22193), .Y(n22370) );
  AOI21XL U6764 ( .A0(n20097), .A1(n20096), .B0(n24849), .Y(n20098) );
  NOR2X1 U6765 ( .A(n22402), .B(n3130), .Y(n22239) );
  OAI2BB1XL U6766 ( .A0N(n25644), .A1N(n25807), .B0(n20965), .Y(n2616) );
  NAND2X1 U6767 ( .A(n22192), .B(n3129), .Y(n22402) );
  AND3X1 U6768 ( .A(n22260), .B(n22395), .C(n22259), .Y(n6168) );
  AOI2BB1XL U6769 ( .A0N(n15714), .A1N(n21000), .B0(n24871), .Y(n15715) );
  OR2X2 U6770 ( .A(n3127), .B(n15767), .Y(n15762) );
  NOR2X1 U6771 ( .A(n3126), .B(n22307), .Y(n22190) );
  AOI21X1 U6772 ( .A0(n23701), .A1(n3229), .B0(n23923), .Y(n23924) );
  NOR2X1 U6773 ( .A(n3126), .B(n22141), .Y(n22197) );
  INVX4 U6774 ( .A(n20473), .Y(n3068) );
  INVX4 U6775 ( .A(n20182), .Y(n3069) );
  CLKINVX3 U6776 ( .A(n15745), .Y(n15808) );
  AOI21XL U6777 ( .A0(n4461), .A1(n3138), .B0(n15923), .Y(n4460) );
  NAND2BX1 U6778 ( .AN(n23603), .B(n3532), .Y(n3531) );
  INVX1 U6779 ( .A(n24606), .Y(n25531) );
  INVX8 U6780 ( .A(n22308), .Y(n3126) );
  INVX4 U6781 ( .A(n8981), .Y(n3071) );
  AOI21XL U6782 ( .A0(n20093), .A1(n20092), .B0(n24717), .Y(n20094) );
  NAND3X1 U6783 ( .A(n5407), .B(n5406), .C(n4714), .Y(n2550) );
  NOR2X1 U6784 ( .A(n9023), .B(n9022), .Y(n9024) );
  CLKINVX3 U6785 ( .A(n8997), .Y(n3073) );
  INVX1 U6786 ( .A(n25556), .Y(n11478) );
  INVXL U6787 ( .A(n20091), .Y(n20093) );
  NAND2X1 U6788 ( .A(n3313), .B(n3312), .Y(n25644) );
  NAND2X1 U6789 ( .A(n4857), .B(n5951), .Y(n2535) );
  AND3XL U6790 ( .A(n5206), .B(n5205), .C(n4711), .Y(n4600) );
  NAND2X1 U6791 ( .A(n3128), .B(n20950), .Y(n3313) );
  NAND2X1 U6792 ( .A(n19104), .B(n20949), .Y(n3312) );
  NAND2X1 U6793 ( .A(n19104), .B(n20950), .Y(n4347) );
  CLKINVX3 U6794 ( .A(n23200), .Y(n3074) );
  NAND2X1 U6795 ( .A(n4976), .B(n25807), .Y(n4975) );
  NAND2X1 U6796 ( .A(n3860), .B(n20353), .Y(n4240) );
  NAND2X1 U6797 ( .A(n3461), .B(n25807), .Y(n3460) );
  NAND2BX1 U6798 ( .AN(n8946), .B(n8945), .Y(n8935) );
  NOR2X1 U6799 ( .A(n25328), .B(n4927), .Y(n24126) );
  BUFX16 U6800 ( .A(n5518), .Y(n3128) );
  NOR2X1 U6801 ( .A(n24170), .B(n25328), .Y(n24173) );
  NOR2X1 U6802 ( .A(n24184), .B(n25328), .Y(n24187) );
  NOR2X1 U6803 ( .A(n24136), .B(n25328), .Y(n24139) );
  AOI21XL U6804 ( .A0(n20089), .A1(n20088), .B0(n20235), .Y(n20090) );
  NOR2X1 U6805 ( .A(n24386), .B(n23778), .Y(n23779) );
  NOR2X1 U6806 ( .A(n4966), .B(n25328), .Y(n24163) );
  NAND2X1 U6807 ( .A(n5011), .B(n20613), .Y(n5002) );
  INVX4 U6808 ( .A(n4950), .Y(n25328) );
  NAND2BX1 U6809 ( .AN(n20076), .B(n20075), .Y(n20064) );
  NAND2X1 U6810 ( .A(n3131), .B(n24123), .Y(n4953) );
  NAND2X1 U6811 ( .A(n24160), .B(n3131), .Y(n3463) );
  NAND2X2 U6812 ( .A(n23751), .B(n3353), .Y(n3998) );
  AND2X2 U6813 ( .A(n20948), .B(n20947), .Y(n20949) );
  INVX1 U6814 ( .A(n20167), .Y(n20168) );
  NAND2BX1 U6815 ( .AN(n15698), .B(n15697), .Y(n15686) );
  AOI21X1 U6816 ( .A0(n3005), .A1(n24051), .B0(n3004), .Y(n3970) );
  CLKINVX3 U6817 ( .A(n23113), .Y(n22461) );
  INVX4 U6818 ( .A(n22281), .Y(n3079) );
  NAND2X1 U6819 ( .A(n20105), .B(n20103), .Y(n20076) );
  OR2X2 U6820 ( .A(n23113), .B(n22124), .Y(n22398) );
  XOR2X1 U6821 ( .A(n8923), .B(n8922), .Y(n20411) );
  XOR2X1 U6822 ( .A(n8933), .B(n8932), .Y(n20432) );
  XNOR2X1 U6823 ( .A(n15480), .B(n15479), .Y(n15872) );
  INVX4 U6824 ( .A(n22124), .Y(n3082) );
  INVX1 U6825 ( .A(n5977), .Y(n4061) );
  XOR2X1 U6826 ( .A(n20052), .B(n20051), .Y(n20188) );
  NAND2X1 U6827 ( .A(n15720), .B(n15718), .Y(n15698) );
  NOR2X1 U6828 ( .A(n20177), .B(n20199), .Y(n20105) );
  AOI21X1 U6829 ( .A0(n8930), .A1(n8762), .B0(n8761), .Y(n8767) );
  XNOR2X1 U6830 ( .A(n15637), .B(n15636), .Y(n25007) );
  XNOR2X1 U6831 ( .A(n8930), .B(n8916), .Y(n20436) );
  AOI21X2 U6832 ( .A0(n8784), .A1(n8783), .B0(n8782), .Y(n8882) );
  NOR2X2 U6833 ( .A(n3321), .B(n3319), .Y(n3234) );
  INVXL U6834 ( .A(n5720), .Y(n5710) );
  NOR2X1 U6835 ( .A(n23604), .B(n4584), .Y(n4821) );
  NAND2X1 U6836 ( .A(n3139), .B(n23539), .Y(n3575) );
  NAND2X1 U6837 ( .A(n3895), .B(n21018), .Y(n21021) );
  INVX1 U6838 ( .A(n9016), .Y(n8953) );
  NOR2X1 U6839 ( .A(n20203), .B(n20204), .Y(n20103) );
  AOI21X2 U6840 ( .A0(n19913), .A1(n19912), .B0(n19911), .Y(n20011) );
  NAND2X1 U6841 ( .A(n3139), .B(n23894), .Y(n3492) );
  INVX1 U6842 ( .A(n8758), .Y(n8930) );
  NOR2BX1 U6843 ( .AN(n15825), .B(n15823), .Y(n15720) );
  XOR2X1 U6844 ( .A(n8910), .B(n8909), .Y(n9015) );
  XNOR2X1 U6845 ( .A(n15680), .B(n15666), .Y(n15820) );
  CLKINVX3 U6846 ( .A(n4508), .Y(n3140) );
  INVX2 U6847 ( .A(n10711), .Y(n5741) );
  NAND2BX1 U6848 ( .AN(n22134), .B(n22133), .Y(n22122) );
  AOI21X1 U6849 ( .A0(n8651), .A1(n8917), .B0(n8650), .Y(n8652) );
  AOI2BB1XL U6850 ( .A0N(n15705), .A1N(n15836), .B0(n15835), .Y(n15706) );
  AOI21X2 U6851 ( .A0(n15533), .A1(n15532), .B0(n15531), .Y(n15632) );
  CLKINVX3 U6852 ( .A(n23431), .Y(n3141) );
  NOR3X1 U6853 ( .A(n22296), .B(n22297), .C(n22157), .Y(n22133) );
  INVXL U6854 ( .A(n20018), .Y(n20033) );
  NAND3X2 U6855 ( .A(n3806), .B(n5700), .C(n5848), .Y(n5658) );
  NOR2X1 U6856 ( .A(n3143), .B(n4636), .Y(n4473) );
  CLKINVX3 U6857 ( .A(n17480), .Y(n19103) );
  XOR2X1 U6858 ( .A(n5696), .B(n5711), .Y(n5695) );
  OR2XL U6859 ( .A(n24251), .B(n24250), .Y(n24252) );
  NAND2X1 U6860 ( .A(n17437), .B(n17433), .Y(n3393) );
  NAND2X1 U6861 ( .A(n8912), .B(n8403), .Y(n8645) );
  AOI21XL U6862 ( .A0(n20071), .A1(n20069), .B0(n20035), .Y(n20039) );
  AOI21X1 U6863 ( .A0(n15382), .A1(n15640), .B0(n15381), .Y(n15507) );
  OR2X1 U6864 ( .A(n22292), .B(n22295), .Y(n22157) );
  NAND2X1 U6865 ( .A(n22155), .B(n22153), .Y(n22134) );
  BUFX2 U6866 ( .A(n6074), .Y(n5740) );
  INVX1 U6867 ( .A(n23495), .Y(n23496) );
  NAND3X1 U6868 ( .A(n6074), .B(n20944), .C(n19073), .Y(n10226) );
  INVX1 U6869 ( .A(n4867), .Y(n3977) );
  BUFX2 U6870 ( .A(n23550), .Y(n5018) );
  NAND2XL U6871 ( .A(n20350), .B(n3357), .Y(n20352) );
  INVX1 U6872 ( .A(n23746), .Y(n5385) );
  INVX1 U6873 ( .A(n20988), .Y(n20989) );
  XOR2X1 U6874 ( .A(n10961), .B(n10960), .Y(n20286) );
  AOI21X1 U6875 ( .A0(n19779), .A1(n20046), .B0(n19778), .Y(n19780) );
  BUFX3 U6876 ( .A(n11464), .Y(n23915) );
  NAND2XL U6877 ( .A(n20927), .B(n20926), .Y(n20928) );
  AOI21X1 U6878 ( .A0(n8461), .A1(n8631), .B0(n8630), .Y(n8890) );
  NAND2X1 U6879 ( .A(n3357), .B(n20738), .Y(n20741) );
  AOI21X1 U6880 ( .A0(n8778), .A1(n8854), .B0(n8777), .Y(n8779) );
  INVX1 U6881 ( .A(n20701), .Y(n23550) );
  XNOR2X1 U6882 ( .A(n15693), .B(n15692), .Y(n15772) );
  CLKINVX3 U6883 ( .A(n23527), .Y(n3146) );
  NAND2X1 U6884 ( .A(n19021), .B(n19019), .Y(n5465) );
  XOR2X1 U6885 ( .A(n22101), .B(n22100), .Y(n22296) );
  XOR2X1 U6886 ( .A(n21956), .B(n21955), .Y(n22244) );
  NOR2X1 U6887 ( .A(n22301), .B(n22302), .Y(n22155) );
  NOR2X1 U6888 ( .A(n22305), .B(n22202), .Y(n22153) );
  NOR2X1 U6889 ( .A(n8637), .B(n8636), .Y(n8924) );
  NOR2X1 U6890 ( .A(n15392), .B(n15674), .Y(n15668) );
  NAND2X1 U6891 ( .A(n3586), .B(n5601), .Y(n20617) );
  CLKINVX3 U6892 ( .A(n4222), .Y(n3084) );
  INVX1 U6893 ( .A(n10963), .Y(n10971) );
  NAND2X1 U6894 ( .A(n20041), .B(n19534), .Y(n19773) );
  NAND2X1 U6895 ( .A(n8637), .B(n8636), .Y(n8926) );
  NAND2XL U6896 ( .A(n3848), .B(n17469), .Y(n5697) );
  AOI21X2 U6897 ( .A0(n21973), .A1(n21972), .B0(n21971), .Y(n22070) );
  XNOR2X1 U6898 ( .A(n22117), .B(n22103), .Y(n22297) );
  NOR2X1 U6899 ( .A(n20923), .B(n20919), .Y(n5394) );
  INVX1 U6900 ( .A(n23456), .Y(n23478) );
  INVX1 U6901 ( .A(n22203), .Y(n22141) );
  NOR2X2 U6902 ( .A(n4142), .B(n23639), .Y(n3862) );
  CLKINVX3 U6903 ( .A(n3931), .Y(n3426) );
  NOR2X2 U6904 ( .A(n5699), .B(n3329), .Y(n3787) );
  CLKINVX3 U6905 ( .A(n20324), .Y(n3344) );
  NOR2X1 U6906 ( .A(n8704), .B(n8703), .Y(n8719) );
  OR2X2 U6907 ( .A(n8629), .B(n8628), .Y(n8461) );
  NAND2XL U6908 ( .A(n8627), .B(n8626), .Y(n8901) );
  INVX1 U6909 ( .A(n13027), .Y(n20672) );
  INVXL U6910 ( .A(n20330), .Y(n20331) );
  NOR2X1 U6911 ( .A(n19765), .B(n19764), .Y(n20053) );
  INVX1 U6912 ( .A(n15621), .Y(n15581) );
  NOR2X1 U6913 ( .A(n15481), .B(n15485), .Y(n15451) );
  INVX1 U6914 ( .A(n23454), .Y(n23455) );
  NOR2X1 U6915 ( .A(n19767), .B(n19766), .Y(n20056) );
  NAND2X1 U6916 ( .A(n13030), .B(n21017), .Y(n4965) );
  NOR2X1 U6917 ( .A(n15384), .B(n15383), .Y(n15674) );
  NOR2X1 U6918 ( .A(n20048), .B(n19892), .Y(n19779) );
  NOR2X1 U6919 ( .A(n8732), .B(n8736), .Y(n8702) );
  NOR2X1 U6920 ( .A(n15589), .B(n15633), .Y(n15569) );
  INVX1 U6921 ( .A(n21017), .Y(n21024) );
  INVX1 U6922 ( .A(n8871), .Y(n8831) );
  NAND2XL U6923 ( .A(n9004), .B(n8823), .Y(n8999) );
  NAND2BX1 U6924 ( .AN(n10653), .B(n10635), .Y(n3326) );
  XNOR2X1 U6925 ( .A(n22129), .B(n22128), .Y(n22203) );
  OR2X2 U6926 ( .A(n19757), .B(n19756), .Y(n19738) );
  NOR2X1 U6927 ( .A(n15447), .B(n15446), .Y(n15481) );
  NAND2XL U6928 ( .A(n15374), .B(n15373), .Y(n15652) );
  NAND2X1 U6929 ( .A(n15571), .B(n15570), .Y(n15621) );
  INVXL U6930 ( .A(n17467), .Y(n20351) );
  AOI21X1 U6931 ( .A0(n11353), .A1(n10952), .B0(n10951), .Y(n10972) );
  INVX2 U6932 ( .A(n20340), .Y(n5717) );
  NOR2X1 U6933 ( .A(n8698), .B(n8697), .Y(n8732) );
  INVXL U6934 ( .A(n10647), .Y(n10634) );
  INVX1 U6935 ( .A(n8839), .Y(n8878) );
  NOR2X1 U6936 ( .A(n19777), .B(n19776), .Y(n19892) );
  AOI21X1 U6937 ( .A0(n21836), .A1(n22104), .B0(n21835), .Y(n21837) );
  OR2XL U6938 ( .A(n24259), .B(n24260), .Y(n24261) );
  XOR2X2 U6939 ( .A(n3805), .B(n4683), .Y(n17463) );
  OR2X1 U6940 ( .A(n8614), .B(n8375), .Y(n8377) );
  OR2X1 U6941 ( .A(n8471), .B(n8614), .Y(n8473) );
  INVX1 U6942 ( .A(n23588), .Y(n20676) );
  INVX1 U6943 ( .A(n18973), .Y(n6091) );
  XOR2X2 U6944 ( .A(n4407), .B(n18922), .Y(n23454) );
  NOR2X1 U6945 ( .A(n15386), .B(n15385), .Y(n15677) );
  NOR2X1 U6946 ( .A(n19833), .B(n19832), .Y(n19848) );
  NOR2X1 U6947 ( .A(n8839), .B(n8883), .Y(n8819) );
  NAND2X1 U6948 ( .A(n8821), .B(n8820), .Y(n8871) );
  NOR2BX1 U6949 ( .AN(n11461), .B(n11458), .Y(n11463) );
  CLKINVX3 U6950 ( .A(n20855), .Y(n3535) );
  NOR2X1 U6951 ( .A(n21830), .B(n22111), .Y(n22105) );
  NOR2X1 U6952 ( .A(n19823), .B(n19822), .Y(n19883) );
  NAND2X2 U6953 ( .A(n10480), .B(n10503), .Y(n4365) );
  XOR2X1 U6954 ( .A(n19686), .B(n3215), .Y(n20145) );
  NOR2X2 U6955 ( .A(n3526), .B(n3527), .Y(n3525) );
  NAND2XL U6956 ( .A(n10503), .B(n10505), .Y(n5220) );
  NOR2X1 U6957 ( .A(n19968), .B(n20012), .Y(n19948) );
  NOR2X1 U6958 ( .A(n19861), .B(n19865), .Y(n19831) );
  CLKBUFX2 U6959 ( .A(n20755), .Y(n20756) );
  OR2X1 U6960 ( .A(n19548), .B(n19748), .Y(n19550) );
  INVX1 U6961 ( .A(n20000), .Y(n19960) );
  INVXL U6962 ( .A(n17445), .Y(n17446) );
  INVX1 U6963 ( .A(n17455), .Y(n20736) );
  NAND2X1 U6964 ( .A(n19940), .B(n19939), .Y(n19977) );
  NOR2X1 U6965 ( .A(n8815), .B(n8814), .Y(n8839) );
  NAND2X1 U6966 ( .A(n8815), .B(n8814), .Y(n8876) );
  NAND3X1 U6967 ( .A(n3809), .B(n3786), .C(n17310), .Y(n3805) );
  XOR2X2 U6968 ( .A(n14638), .B(n14477), .Y(n14663) );
  NAND2X1 U6969 ( .A(n8817), .B(n8816), .Y(n8884) );
  INVX1 U6970 ( .A(n10729), .Y(n5097) );
  AOI21XL U6971 ( .A0(n15347), .A1(n15346), .B0(n15345), .Y(n15348) );
  INVX1 U6972 ( .A(n10197), .Y(n10199) );
  INVX1 U6973 ( .A(n12814), .Y(n12811) );
  NOR2X1 U6974 ( .A(n19827), .B(n19826), .Y(n19861) );
  OR2X1 U6975 ( .A(n19749), .B(n19748), .Y(n19751) );
  NOR2X1 U6976 ( .A(n21822), .B(n21821), .Y(n22111) );
  NAND2X1 U6977 ( .A(n19950), .B(n19949), .Y(n20000) );
  INVX1 U6978 ( .A(n12845), .Y(n12847) );
  INVX1 U6979 ( .A(n20282), .Y(n20280) );
  INVX1 U6980 ( .A(n14552), .Y(n14567) );
  NAND2X1 U6981 ( .A(n5272), .B(n14636), .Y(n14477) );
  NOR2X1 U6982 ( .A(n8503), .B(n3154), .Y(n8769) );
  NAND2BX1 U6983 ( .AN(n17296), .B(n4151), .Y(n4150) );
  NOR2X1 U6984 ( .A(n8661), .B(n3154), .Y(n8790) );
  NAND2X2 U6985 ( .A(n5059), .B(n17373), .Y(n17381) );
  NAND2X2 U6986 ( .A(n3951), .B(n17351), .Y(n17356) );
  XOR2X2 U6987 ( .A(n3588), .B(n7432), .Y(n10741) );
  NAND2XL U6988 ( .A(n21740), .B(n3222), .Y(n22186) );
  INVX1 U6989 ( .A(n20853), .Y(n20866) );
  INVX1 U6990 ( .A(n20869), .Y(n20870) );
  INVX1 U6991 ( .A(n20759), .Y(n20845) );
  AND2X1 U6992 ( .A(n8610), .B(n8822), .Y(n8398) );
  NOR2X1 U6993 ( .A(n8511), .B(n3154), .Y(n8805) );
  NAND2BX2 U6994 ( .AN(n20637), .B(n9198), .Y(n20642) );
  AOI21X1 U6995 ( .A0(n10948), .A1(n10983), .B0(n10947), .Y(n11393) );
  AOI21XL U6996 ( .A0(n10651), .A1(n10650), .B0(n10649), .Y(n10652) );
  NAND2X1 U6997 ( .A(n5667), .B(n17352), .Y(n3951) );
  AND2X2 U6998 ( .A(n17341), .B(n17344), .Y(n17347) );
  INVX1 U6999 ( .A(n14637), .Y(n5272) );
  NAND2X1 U7000 ( .A(n14611), .B(n14610), .Y(n14612) );
  NAND2X1 U7001 ( .A(n14570), .B(n14569), .Y(n14571) );
  AND2X2 U7002 ( .A(n10058), .B(n10057), .Y(n3241) );
  NAND2X1 U7003 ( .A(n8295), .B(n8795), .Y(n8797) );
  AOI2BB2X1 U7004 ( .B0(n8550), .B1(n3157), .A0N(n3157), .A1N(n8453), .Y(n8661) );
  NOR2X1 U7005 ( .A(n21921), .B(n21925), .Y(n21891) );
  AOI2BB2X1 U7006 ( .B0(n8345), .B1(n3157), .A0N(n3157), .A1N(n8406), .Y(n8503) );
  NOR2X1 U7007 ( .A(n21824), .B(n21823), .Y(n22114) );
  AOI2BB2XL U7008 ( .B0(n8452), .B1(n3157), .A0N(n3157), .A1N(n8451), .Y(n8662) );
  AND2X1 U7009 ( .A(n15355), .B(n15572), .Y(n15147) );
  NAND2X1 U7010 ( .A(n4360), .B(n3150), .Y(n10505) );
  INVX1 U7011 ( .A(n22059), .Y(n22019) );
  NOR2X1 U7012 ( .A(n22027), .B(n22071), .Y(n22008) );
  AOI21X1 U7013 ( .A0(n12835), .A1(n12853), .B0(n12852), .Y(n12854) );
  NOR2X1 U7014 ( .A(n8570), .B(n8669), .Y(n8795) );
  NAND2X1 U7015 ( .A(n22010), .B(n22009), .Y(n22059) );
  INVX1 U7016 ( .A(n15359), .Y(n15256) );
  NOR2X1 U7017 ( .A(n21893), .B(n21892), .Y(n21908) );
  NAND2X1 U7018 ( .A(n19424), .B(n19929), .Y(n19931) );
  NOR2X1 U7019 ( .A(n19789), .B(n19807), .Y(n19919) );
  NOR2X1 U7020 ( .A(n21885), .B(n21884), .Y(n21938) );
  NAND2X1 U7021 ( .A(n22000), .B(n21999), .Y(n22036) );
  NAND2X1 U7022 ( .A(n10177), .B(n10464), .Y(n10178) );
  NAND2X1 U7023 ( .A(n18408), .B(n18407), .Y(n18914) );
  NOR2X1 U7024 ( .A(n8603), .B(n3154), .Y(n8822) );
  AOI2BB1X2 U7025 ( .A0N(n12836), .A1N(n4056), .B0(n4036), .Y(n4035) );
  XNOR2X1 U7026 ( .A(n3570), .B(n7368), .Y(n3569) );
  INVXL U7027 ( .A(n17371), .Y(n3149) );
  NOR2X1 U7028 ( .A(n8570), .B(n8676), .Y(n8800) );
  INVX1 U7029 ( .A(n10468), .Y(n3306) );
  INVX1 U7030 ( .A(n18999), .Y(n19002) );
  NOR2X4 U7031 ( .A(n15359), .B(n15355), .Y(n15046) );
  NAND2X1 U7032 ( .A(n19424), .B(n19924), .Y(n19926) );
  AND2X2 U7033 ( .A(n12858), .B(n12979), .Y(n4615) );
  AOI2BB2XL U7034 ( .B0(n15424), .B1(n3016), .A0N(n3016), .A1N(n15153), .Y(
        n15244) );
  AOI2BB2XL U7035 ( .B0(n15416), .B1(n3016), .A0N(n3016), .A1N(n15210), .Y(
        n15224) );
  NAND2X2 U7036 ( .A(n15329), .B(n15040), .Y(n15359) );
  AOI2BB2XL U7037 ( .B0(n6194), .B1(n15182), .A0N(n3156), .A1N(n15181), .Y(
        n15402) );
  AOI2BB2XL U7038 ( .B0(n15199), .B1(n3016), .A0N(n3016), .A1N(n15198), .Y(
        n15409) );
  NOR2X1 U7039 ( .A(n19739), .B(n19797), .Y(n19924) );
  AND2X2 U7040 ( .A(n17209), .B(n17208), .Y(n4588) );
  NOR2X1 U7041 ( .A(n19739), .B(n19804), .Y(n19929) );
  AND3X1 U7042 ( .A(n21670), .B(n21669), .C(n21859), .Y(n4623) );
  AOI21X1 U7043 ( .A0(n12883), .A1(n12926), .B0(n12882), .Y(n12884) );
  AOI2BB2X1 U7044 ( .B0(n19729), .B1(n19542), .A0N(n19542), .A1N(n19728), .Y(
        n19789) );
  AOI21X1 U7045 ( .A0(n19011), .A1(n19010), .B0(n19009), .Y(n19012) );
  AOI21X1 U7046 ( .A0(n7364), .A1(n7363), .B0(n7362), .Y(n3570) );
  INVX1 U7047 ( .A(n17418), .Y(n3628) );
  INVX1 U7048 ( .A(n18963), .Y(n18957) );
  AOI21X1 U7049 ( .A0(n18948), .A1(n18947), .B0(n18946), .Y(n18949) );
  AND2X2 U7050 ( .A(n15416), .B(n15336), .Y(n15544) );
  NAND2X1 U7051 ( .A(n8601), .B(n8434), .Y(n8570) );
  NAND3X1 U7052 ( .A(n7437), .B(n7442), .C(n7443), .Y(n5128) );
  NOR4BXL U7053 ( .AN(n21736), .B(n21735), .C(n21734), .D(n21733), .Y(n21738)
         );
  INVX1 U7054 ( .A(n20641), .Y(n20647) );
  NAND2X2 U7055 ( .A(n12863), .B(n12858), .Y(n12833) );
  AND2X1 U7056 ( .A(n19730), .B(n19951), .Y(n19529) );
  NAND2X1 U7057 ( .A(n10574), .B(n10562), .Y(n10585) );
  AOI2BB2XL U7058 ( .B0(n15119), .B1(n3016), .A0N(n3016), .A1N(n15181), .Y(
        n15263) );
  NOR3XL U7059 ( .A(n21695), .B(n21694), .C(n21693), .Y(n21739) );
  INVX1 U7060 ( .A(n17230), .Y(n17211) );
  ADDFHX2 U7061 ( .A(n9372), .B(n9371), .CI(n9370), .CO(n10132), .S(n10131) );
  INVX1 U7062 ( .A(n23662), .Y(n23659) );
  NAND2X1 U7063 ( .A(n4619), .B(n10607), .Y(n4589) );
  NOR2X1 U7064 ( .A(n17415), .B(n17417), .Y(n17294) );
  NAND2X1 U7065 ( .A(n3036), .B(n19714), .Y(n19600) );
  INVX1 U7066 ( .A(n24034), .Y(n14692) );
  OR2X2 U7067 ( .A(n20640), .B(n20639), .Y(n20641) );
  INVX1 U7068 ( .A(n10614), .Y(n10631) );
  NOR2X4 U7069 ( .A(n19748), .B(n19730), .Y(n19424) );
  AOI2BB2XL U7070 ( .B0(n15184), .B1(n3016), .A0N(n3016), .A1N(n15183), .Y(
        n15401) );
  NAND2X1 U7071 ( .A(n18900), .B(n18899), .Y(n18901) );
  NAND2X1 U7072 ( .A(n3156), .B(n15184), .Y(n15262) );
  OAI21X2 U7073 ( .A0(n5380), .A1(n3008), .B0(n5378), .Y(n10123) );
  AND2X2 U7074 ( .A(n17328), .B(n17313), .Y(n4604) );
  NAND2X1 U7075 ( .A(n3153), .B(n12895), .Y(n12878) );
  OR2XL U7076 ( .A(n18841), .B(n18843), .Y(n4675) );
  CLKINVX3 U7077 ( .A(n3157), .Y(n3087) );
  NAND2XL U7078 ( .A(n21506), .B(n22011), .Y(n22013) );
  BUFX3 U7079 ( .A(n3423), .Y(n3422) );
  NAND2BX1 U7080 ( .AN(n10500), .B(n10555), .Y(n10556) );
  NAND2X1 U7081 ( .A(n12924), .B(n12923), .Y(n4664) );
  INVX1 U7082 ( .A(n12896), .Y(n3153) );
  AND2X2 U7083 ( .A(n10638), .B(n10637), .Y(n4628) );
  ADDFHX1 U7084 ( .A(n14138), .B(n14137), .CI(n14136), .CO(n14320), .S(n14317)
         );
  AND2X2 U7085 ( .A(n8598), .B(n9027), .Y(n8668) );
  CLKINVX3 U7086 ( .A(n3016), .Y(n3156) );
  INVX1 U7087 ( .A(n9268), .Y(n5077) );
  NAND2X2 U7088 ( .A(n17236), .B(n16866), .Y(n3366) );
  AND2X2 U7089 ( .A(n10641), .B(n10551), .Y(n4665) );
  XOR2X1 U7090 ( .A(n9764), .B(n3280), .Y(n3279) );
  INVX2 U7091 ( .A(n4591), .Y(n8606) );
  NAND2X2 U7092 ( .A(n17328), .B(n17331), .Y(n3328) );
  INVX1 U7093 ( .A(n18886), .Y(n18900) );
  NAND2X1 U7094 ( .A(n18863), .B(n18862), .Y(n18864) );
  AOI22XL U7095 ( .A0(n21659), .A1(n3037), .B0(n3171), .B1(n21658), .Y(n21872)
         );
  NAND2XL U7096 ( .A(n10290), .B(n10291), .Y(n5527) );
  AOI22X1 U7097 ( .A0(n3167), .A1(n15132), .B0(n3038), .B1(n15055), .Y(n15424)
         );
  AOI22X1 U7098 ( .A0(n3167), .A1(n15112), .B0(n15120), .B1(n15055), .Y(n15416) );
  ADDFHX1 U7099 ( .A(n14068), .B(n14067), .CI(n14066), .CO(n14161), .S(n14037)
         );
  NAND2BX2 U7100 ( .AN(n10039), .B(n3238), .Y(n3253) );
  NAND2BX1 U7101 ( .AN(n24033), .B(n24029), .Y(n24030) );
  ADDFHX1 U7102 ( .A(n13829), .B(n13828), .CI(n13827), .CO(n13907), .S(n13830)
         );
  ADDFHX2 U7103 ( .A(n16154), .B(n16153), .CI(n16152), .CO(n16854), .S(n16853)
         );
  NAND2X2 U7104 ( .A(n23955), .B(n15345), .Y(n15363) );
  NAND2X1 U7105 ( .A(n18992), .B(n18997), .Y(n18716) );
  CLKINVX3 U7106 ( .A(n7423), .Y(n7442) );
  NOR2X1 U7107 ( .A(n15055), .B(n15120), .Y(n15184) );
  NOR2XL U7108 ( .A(n21641), .B(n3171), .Y(n21958) );
  NAND2X1 U7109 ( .A(n6113), .B(n4932), .Y(n12768) );
  AND2X2 U7110 ( .A(n10584), .B(n10583), .Y(n4681) );
  INVX1 U7111 ( .A(n10500), .Y(n10641) );
  INVXL U7112 ( .A(n13753), .Y(n5292) );
  NOR2XL U7113 ( .A(n21618), .B(n3171), .Y(n21898) );
  INVX1 U7114 ( .A(n12906), .Y(n12893) );
  INVX1 U7115 ( .A(n17227), .Y(n17297) );
  INVX1 U7116 ( .A(n17314), .Y(n4942) );
  NOR2X4 U7117 ( .A(n21787), .B(n21803), .Y(n21506) );
  OR2X2 U7118 ( .A(n9192), .B(n10670), .Y(n9191) );
  AND2X2 U7119 ( .A(n3000), .B(n18931), .Y(n4608) );
  NAND2X1 U7120 ( .A(n4981), .B(n6002), .Y(n4376) );
  OAI2BB1X1 U7121 ( .A0N(n10063), .A1N(n10064), .B0(n3262), .Y(n9416) );
  NAND2X1 U7122 ( .A(n8225), .B(n8268), .Y(n8226) );
  NOR2X1 U7123 ( .A(n10575), .B(n10582), .Y(n10562) );
  AOI21X1 U7124 ( .A0(n7819), .A1(n7818), .B0(n7817), .Y(n7820) );
  AND2X2 U7125 ( .A(n7325), .B(n7320), .Y(n7311) );
  AND2X2 U7126 ( .A(n21864), .B(n21793), .Y(n21989) );
  CLKINVX3 U7127 ( .A(n19457), .Y(n3166) );
  NAND2X1 U7128 ( .A(n14495), .B(n14490), .Y(n14491) );
  AND2X2 U7129 ( .A(n19683), .B(n3215), .Y(n19796) );
  ADDFHX1 U7130 ( .A(n10394), .B(n10393), .CI(n10392), .CO(n10476), .S(n10473)
         );
  NOR2X1 U7131 ( .A(n10502), .B(n10501), .Y(n10500) );
  XOR2X1 U7132 ( .A(n9414), .B(n9415), .Y(n5309) );
  NAND2X1 U7133 ( .A(n10481), .B(n10482), .Y(n10637) );
  NOR2X1 U7134 ( .A(n21658), .B(n3171), .Y(n21994) );
  NAND2X1 U7135 ( .A(n8286), .B(n8276), .Y(n8277) );
  INVX1 U7136 ( .A(n9192), .Y(n20639) );
  NAND2X2 U7137 ( .A(n5477), .B(n5476), .Y(n17646) );
  OR2XL U7138 ( .A(n23960), .B(n23167), .Y(n23172) );
  ADDFHX2 U7139 ( .A(n13759), .B(n13758), .CI(n13757), .CO(n13826), .S(n13760)
         );
  XOR3X2 U7140 ( .A(n10318), .B(n10316), .C(n10317), .Y(n10290) );
  NAND2X1 U7141 ( .A(n12794), .B(n12807), .Y(n12824) );
  AOI21X1 U7142 ( .A0(n8273), .A1(n8272), .B0(n8271), .Y(n8294) );
  NAND2X2 U7143 ( .A(n3611), .B(n3610), .Y(n3609) );
  INVX1 U7144 ( .A(n8279), .Y(n8286) );
  XOR2X2 U7145 ( .A(n19423), .B(n19422), .Y(n19730) );
  NAND2X1 U7146 ( .A(n18979), .B(n18709), .Y(n19006) );
  XNOR2X1 U7147 ( .A(n9830), .B(n9831), .Y(n5177) );
  INVX1 U7148 ( .A(n16776), .Y(n3615) );
  AND2X2 U7149 ( .A(n10680), .B(n9139), .Y(n9192) );
  OAI21XL U7150 ( .A0(n19382), .A1(n19396), .B0(n19398), .Y(n19357) );
  NAND2X1 U7151 ( .A(n7449), .B(n7448), .Y(n7450) );
  NAND2X1 U7152 ( .A(n4689), .B(n10723), .Y(n10724) );
  NOR2X1 U7153 ( .A(n10558), .B(n10557), .Y(n10575) );
  OAI2BB1XL U7154 ( .A0N(n14084), .A1N(n4276), .B0(n4274), .Y(n14108) );
  NOR2X1 U7155 ( .A(n3039), .B(n19642), .Y(n19502) );
  NOR2X1 U7156 ( .A(n3038), .B(n15315), .Y(n15120) );
  NAND2X1 U7157 ( .A(n12840), .B(n12849), .Y(n12850) );
  NAND2X1 U7158 ( .A(n7306), .B(n7489), .Y(n7307) );
  NOR2X1 U7159 ( .A(n9139), .B(n10680), .Y(n10670) );
  ADDFHX1 U7160 ( .A(n10016), .B(n10015), .CI(n10014), .CO(n10042), .S(n10036)
         );
  NAND2X1 U7161 ( .A(n3172), .B(n21769), .Y(n21658) );
  AOI21X1 U7162 ( .A0(n10965), .A1(n10954), .B0(n10953), .Y(n11015) );
  AND2X2 U7163 ( .A(n12977), .B(n12976), .Y(n4678) );
  NOR2XL U7164 ( .A(n5992), .B(n12787), .Y(n5991) );
  NOR2X2 U7165 ( .A(n12510), .B(n12509), .Y(n12905) );
  OAI21X1 U7166 ( .A0(n10064), .A1(n10063), .B0(n10062), .Y(n3262) );
  ADDFHX1 U7167 ( .A(n9294), .B(n9293), .CI(n9292), .CO(n9347), .S(n9372) );
  NOR2X1 U7168 ( .A(n14339), .B(n14338), .Y(n14506) );
  OAI21X2 U7169 ( .A0(n3907), .A1(n3906), .B0(n3905), .Y(n12473) );
  OAI21XL U7170 ( .A0(n4458), .A1(n15010), .B0(n15012), .Y(n14973) );
  CLKINVX3 U7171 ( .A(n12112), .Y(n3473) );
  NAND2X1 U7172 ( .A(n14971), .B(n15011), .Y(n14972) );
  NAND2X1 U7173 ( .A(n7431), .B(n7430), .Y(n7432) );
  AND2X1 U7174 ( .A(n10650), .B(n10648), .Y(n4703) );
  NAND2BX1 U7175 ( .AN(n16805), .B(n3683), .Y(n3682) );
  NAND2X1 U7176 ( .A(n23810), .B(n8223), .Y(n8269) );
  AND2X2 U7177 ( .A(n12871), .B(n12870), .Y(n4684) );
  NAND2X1 U7178 ( .A(n23816), .B(n8224), .Y(n8268) );
  ADDFHX2 U7179 ( .A(n16086), .B(n16085), .CI(n16084), .CO(n16079), .S(n16783)
         );
  ADDFHX1 U7180 ( .A(n12671), .B(n12670), .CI(n12669), .CO(n12769), .S(n12767)
         );
  CLKBUFX2 U7181 ( .A(n12940), .Y(n12972) );
  OAI21XL U7182 ( .A0(n17027), .A1(n17028), .B0(n17026), .Y(n5661) );
  XOR2X1 U7183 ( .A(n17027), .B(n17028), .Y(n5664) );
  AND2X2 U7184 ( .A(n17355), .B(n17310), .Y(n4679) );
  INVXL U7185 ( .A(n12667), .Y(n5039) );
  INVXL U7186 ( .A(n12415), .Y(n6002) );
  NAND2X1 U7187 ( .A(n7873), .B(n10726), .Y(n7870) );
  INVX1 U7188 ( .A(n7308), .Y(n7325) );
  OAI22X1 U7189 ( .A0(n16766), .A1(n3946), .B0(n3945), .B1(n3944), .Y(n3943)
         );
  NAND2X1 U7190 ( .A(n3170), .B(n12867), .Y(n4627) );
  ADDFHX1 U7191 ( .A(n13910), .B(n13909), .CI(n13908), .CO(n13946), .S(n13943)
         );
  ADDFHX1 U7192 ( .A(n13239), .B(n13238), .CI(n13237), .CO(n13309), .S(n13240)
         );
  NAND2X1 U7193 ( .A(n19355), .B(n19397), .Y(n19356) );
  INVX1 U7194 ( .A(n16775), .Y(n3614) );
  OAI21XL U7195 ( .A0(n4017), .A1(n4016), .B0(n4015), .Y(n12421) );
  NAND2X1 U7196 ( .A(n19421), .B(n19420), .Y(n19422) );
  INVXL U7197 ( .A(n13752), .Y(n5291) );
  ADDFHX1 U7198 ( .A(n10031), .B(n10030), .CI(n10029), .CO(n10033), .S(n10007)
         );
  OR2XL U7199 ( .A(n23844), .B(n8281), .Y(n8280) );
  NAND2X1 U7200 ( .A(n17355), .B(n4634), .Y(n17133) );
  AND2X2 U7201 ( .A(n18953), .B(n18952), .Y(n18954) );
  ADDFHX1 U7202 ( .A(n10082), .B(n10081), .CI(n10080), .CO(n10102), .S(n10106)
         );
  INVXL U7203 ( .A(n9523), .Y(n5522) );
  AND2X2 U7204 ( .A(n8287), .B(n23690), .Y(n6178) );
  NAND2XL U7205 ( .A(n14994), .B(n15012), .Y(n4459) );
  NAND2X1 U7206 ( .A(n20656), .B(n20655), .Y(n20657) );
  ADDFHX1 U7207 ( .A(n9473), .B(n9472), .CI(n9471), .CO(n9523), .S(n9456) );
  NAND2X1 U7208 ( .A(n7722), .B(n7727), .Y(n7788) );
  ADDFHX2 U7209 ( .A(n10168), .B(n10167), .CI(n10166), .CO(n10293), .S(n10149)
         );
  ADDFHX1 U7210 ( .A(n10153), .B(n10152), .CI(n10151), .CO(n10318), .S(n10173)
         );
  XNOR2X1 U7211 ( .A(n9181), .B(n9180), .Y(n23776) );
  NAND2X1 U7212 ( .A(n7305), .B(n7304), .Y(n7489) );
  OAI21XL U7213 ( .A0(n4357), .A1(n2976), .B0(n10297), .Y(n4355) );
  NAND2X1 U7214 ( .A(n7269), .B(n7268), .Y(n7439) );
  ADDFHX2 U7215 ( .A(n18593), .B(n18592), .CI(n18591), .CO(n18677), .S(n18674)
         );
  XNOR2X1 U7216 ( .A(n5069), .B(n9316), .Y(n5072) );
  INVXL U7217 ( .A(n5069), .Y(n3453) );
  OR2X2 U7218 ( .A(n10572), .B(n10571), .Y(n10650) );
  INVX1 U7219 ( .A(n19409), .Y(n19406) );
  NAND2BX2 U7220 ( .AN(n20649), .B(n18971), .Y(n20655) );
  NAND2X1 U7221 ( .A(n7776), .B(n7775), .Y(n7777) );
  NAND2X1 U7222 ( .A(n7772), .B(n7657), .Y(n7522) );
  XNOR2X1 U7223 ( .A(n11919), .B(n3658), .Y(n11902) );
  INVX1 U7224 ( .A(n23183), .Y(n8223) );
  NAND2BX2 U7225 ( .AN(n17128), .B(n5083), .Y(n17355) );
  XOR2X1 U7226 ( .A(n21449), .B(n21448), .Y(n4618) );
  AND2X2 U7227 ( .A(n18962), .B(n18959), .Y(n4596) );
  NAND2XL U7228 ( .A(n3836), .B(n3835), .Y(n17848) );
  ADDFHX2 U7229 ( .A(n17025), .B(n17024), .CI(n17023), .CO(n17026), .S(n17014)
         );
  ADDFHX1 U7230 ( .A(n13704), .B(n13703), .CI(n13702), .CO(n13744), .S(n13805)
         );
  OAI21X1 U7231 ( .A0(n4429), .A1(n4428), .B0(n4427), .Y(n11766) );
  INVX1 U7232 ( .A(n23181), .Y(n8274) );
  NAND2BX1 U7233 ( .AN(n3966), .B(n11971), .Y(n4998) );
  NOR2X1 U7234 ( .A(n21580), .B(n21572), .Y(n21769) );
  NOR2X1 U7235 ( .A(n4793), .B(n15018), .Y(n15023) );
  NAND2XL U7236 ( .A(n12676), .B(n12677), .Y(n3978) );
  XNOR2X1 U7237 ( .A(n12679), .B(n12680), .Y(n4032) );
  NAND2XL U7238 ( .A(n3778), .B(n16818), .Y(n3777) );
  NAND3X1 U7239 ( .A(n4787), .B(n4793), .C(n24020), .Y(n14924) );
  ADDFHX1 U7240 ( .A(n18574), .B(n18573), .CI(n18572), .CO(n18684), .S(n18681)
         );
  NAND2X1 U7241 ( .A(n4787), .B(n14970), .Y(n15011) );
  INVXL U7242 ( .A(n12680), .Y(n4905) );
  AND2X2 U7243 ( .A(n12817), .B(n12815), .Y(n4686) );
  NAND2BXL U7244 ( .AN(n14084), .B(n4278), .Y(n4275) );
  ADDFHX1 U7245 ( .A(n13856), .B(n13855), .CI(n13854), .CO(n13903), .S(n13827)
         );
  OAI2BB1X1 U7246 ( .A0N(n16829), .A1N(n16828), .B0(n3774), .Y(n16821) );
  AND2X2 U7247 ( .A(n19416), .B(n24300), .Y(n6200) );
  NAND2X1 U7248 ( .A(n24433), .B(n19411), .Y(n19415) );
  OR2XL U7249 ( .A(n24433), .B(n19411), .Y(n19410) );
  ADDFHX1 U7250 ( .A(n13850), .B(n13849), .CI(n13848), .CO(n13868), .S(n13856)
         );
  OR2XL U7251 ( .A(M6_mult_x_15_n647), .B(M6_mult_x_15_n656), .Y(n10927) );
  OR2XL U7252 ( .A(M6_mult_x_15_n438), .B(M6_mult_x_15_n441), .Y(n11011) );
  XNOR2X1 U7253 ( .A(n20651), .B(n4522), .Y(n20649) );
  ADDFHX1 U7254 ( .A(n13894), .B(n13893), .CI(n13892), .CO(n13921), .S(n13881)
         );
  AND2X2 U7255 ( .A(n10665), .B(n10664), .Y(n4701) );
  NOR2X1 U7256 ( .A(n24341), .B(n19353), .Y(n19396) );
  NAND2X1 U7257 ( .A(n24341), .B(n19353), .Y(n19398) );
  ADDFHX1 U7258 ( .A(n9263), .B(n9262), .CI(n9261), .CO(n9284), .S(n9313) );
  INVXL U7259 ( .A(n11825), .Y(n4026) );
  XNOR2X2 U7260 ( .A(n5244), .B(n5073), .Y(n5069) );
  NAND2X1 U7261 ( .A(n24092), .B(n19352), .Y(n19359) );
  NOR2XL U7262 ( .A(n16763), .B(n16762), .Y(n3788) );
  ADDFHX1 U7263 ( .A(n9308), .B(n9307), .CI(n9306), .CO(n9316), .S(n9390) );
  INVXL U7264 ( .A(n16764), .Y(n3944) );
  NOR2X1 U7265 ( .A(n24295), .B(n19403), .Y(n19419) );
  NAND2X1 U7266 ( .A(n24295), .B(n19403), .Y(n19420) );
  ADDFHX1 U7267 ( .A(n13796), .B(n13795), .CI(n13794), .CO(n13855), .S(n13782)
         );
  XNOR2X1 U7268 ( .A(n12133), .B(n3387), .Y(n12135) );
  NAND2X1 U7269 ( .A(n9149), .B(n10678), .Y(n9145) );
  NAND2X1 U7270 ( .A(n24072), .B(n19354), .Y(n19397) );
  OAI21XL U7271 ( .A0(n8161), .A1(n8198), .B0(n8197), .Y(n23185) );
  AND2X2 U7272 ( .A(n17380), .B(n17378), .Y(n4682) );
  OR2X2 U7273 ( .A(n23640), .B(n23639), .Y(n5739) );
  AND4X2 U7274 ( .A(n19344), .B(n19343), .C(n19342), .D(n19341), .Y(n19345) );
  NOR2XL U7275 ( .A(n11972), .B(n11973), .Y(n3966) );
  INVXL U7276 ( .A(n11972), .Y(n4999) );
  XOR2X2 U7277 ( .A(n21505), .B(n21504), .Y(n21803) );
  NOR2X1 U7278 ( .A(n18980), .B(n18988), .Y(n18709) );
  INVXL U7279 ( .A(n11973), .Y(n5000) );
  OAI2BB1X1 U7280 ( .A0N(n17002), .A1N(n17001), .B0(n5950), .Y(n17013) );
  INVX4 U7281 ( .A(n21560), .Y(n3096) );
  AND2X2 U7282 ( .A(n7744), .B(n7745), .Y(n4610) );
  OAI22X1 U7283 ( .A0(n8799), .A1(n3017), .B0(n3040), .B1(n8798), .Y(n8814) );
  NOR2X1 U7284 ( .A(n17126), .B(n17125), .Y(n17309) );
  OAI21XL U7285 ( .A0(n17796), .A1(n17797), .B0(n17795), .Y(n5927) );
  ADDFHX1 U7286 ( .A(n17019), .B(n17018), .CI(n17017), .CO(n17028), .S(n17023)
         );
  OAI21X1 U7287 ( .A0(n18360), .A1(n18361), .B0(n18359), .Y(n4090) );
  AND2X2 U7288 ( .A(n15038), .B(n24020), .Y(n6195) );
  NOR2BX1 U7289 ( .AN(n7869), .B(n7868), .Y(n7877) );
  ADDFHX1 U7290 ( .A(n17815), .B(n17814), .CI(n17813), .CO(n18581), .S(n17816)
         );
  OAI22XL U7291 ( .A0(n18295), .A1(n18294), .B0(n5422), .B1(n5421), .Y(n18296)
         );
  OR2XL U7292 ( .A(n9931), .B(n9930), .Y(n9929) );
  ADDFHX1 U7293 ( .A(n12610), .B(n12609), .CI(n12608), .CO(n12775), .S(n12772)
         );
  ADDFHX1 U7294 ( .A(n9611), .B(n9610), .CI(n9609), .CO(n10078), .S(n9649) );
  NAND2XL U7295 ( .A(n17128), .B(n17127), .Y(n17310) );
  AND2X2 U7296 ( .A(n18966), .B(n18967), .Y(n4685) );
  OR2XL U7297 ( .A(n13111), .B(n13110), .Y(n13109) );
  OAI22X1 U7298 ( .A0(n8794), .A1(n3017), .B0(n3040), .B1(n8793), .Y(n8812) );
  NAND2XL U7299 ( .A(n17643), .B(n17644), .Y(n3835) );
  ADDFHX2 U7300 ( .A(n11736), .B(n11735), .CI(n11734), .CO(n11752), .S(n11824)
         );
  NOR2X1 U7301 ( .A(n7681), .B(n7746), .Y(n7722) );
  NAND2X1 U7302 ( .A(n3040), .B(n8180), .Y(n8166) );
  NAND2X1 U7303 ( .A(n3040), .B(n8199), .Y(n8172) );
  OAI21XL U7304 ( .A0(n13738), .A1(n14227), .B0(n4670), .Y(n13733) );
  OAI21XL U7305 ( .A0(n10458), .A1(n3174), .B0(n5752), .Y(n10455) );
  OR4XL U7306 ( .A(n24390), .B(n24300), .C(n24433), .D(n24309), .Y(n20136) );
  INVXL U7307 ( .A(n12679), .Y(n4904) );
  NAND2X1 U7308 ( .A(n8482), .B(n8207), .Y(n8168) );
  NAND2X1 U7309 ( .A(n3040), .B(n8203), .Y(n8170) );
  ADDFHX1 U7310 ( .A(n11970), .B(n11969), .CI(n11968), .CO(n12674), .S(n11971)
         );
  ADDFHX2 U7311 ( .A(n11804), .B(n11803), .CI(n11802), .CO(n11825), .S(n11859)
         );
  NAND2X1 U7312 ( .A(n7483), .B(n7482), .Y(n7488) );
  AOI2BB1X1 U7313 ( .A0N(n23645), .A1N(n21170), .B0(n21169), .Y(mul5_out[31])
         );
  INVX1 U7314 ( .A(n17378), .Y(n17379) );
  NAND2X1 U7315 ( .A(n21503), .B(n21502), .Y(n21504) );
  NAND2X1 U7316 ( .A(n7807), .B(n7749), .Y(n7750) );
  AND2XL U7317 ( .A(n6667), .B(n6666), .Y(n6671) );
  NOR2X1 U7318 ( .A(n21643), .B(n21709), .Y(n21572) );
  ADDFHX1 U7319 ( .A(n13675), .B(n13674), .CI(n13673), .CO(n13740), .S(n13703)
         );
  ADDFHX1 U7320 ( .A(n11942), .B(n11941), .CI(n11940), .CO(n11973), .S(n11939)
         );
  ADDFHX1 U7321 ( .A(n11739), .B(n11738), .CI(n11737), .CO(n11734), .S(n11828)
         );
  NOR2X1 U7322 ( .A(n12790), .B(n12789), .Y(n12812) );
  OAI21X1 U7323 ( .A0(n3287), .A1(n9651), .B0(n3294), .Y(n9646) );
  NOR2X1 U7324 ( .A(n18705), .B(n18704), .Y(n18980) );
  INVXL U7325 ( .A(n3814), .Y(n3813) );
  INVXL U7326 ( .A(n17844), .Y(n5903) );
  INVXL U7327 ( .A(n17843), .Y(n5902) );
  NOR2X1 U7328 ( .A(n17376), .B(n17383), .Y(n17139) );
  XNOR2X1 U7329 ( .A(n9377), .B(n3269), .Y(n3268) );
  NAND2X1 U7330 ( .A(n17141), .B(n17140), .Y(n17392) );
  ADDFHX1 U7331 ( .A(n18474), .B(n18473), .CI(n18472), .CO(n18688), .S(n18685)
         );
  OR2XL U7332 ( .A(n9910), .B(n9909), .Y(n9908) );
  NAND4X1 U7333 ( .A(n24433), .B(n24092), .C(n24341), .D(n24295), .Y(n19308)
         );
  INVX1 U7334 ( .A(n16046), .Y(n4154) );
  AOI2BB2X2 U7335 ( .B0(n23637), .B1(n23638), .A0N(n23638), .A1N(n23637), .Y(
        n23634) );
  XOR2X1 U7336 ( .A(n12175), .B(n4005), .Y(n4881) );
  ADDFHX2 U7337 ( .A(n18571), .B(n18570), .CI(n18569), .CO(n18575), .S(n18595)
         );
  ADDFHX2 U7338 ( .A(n16811), .B(n16810), .CI(n16809), .CO(n16803), .S(n16826)
         );
  XOR2X1 U7339 ( .A(n9246), .B(n4311), .Y(n4310) );
  ADDFHX2 U7340 ( .A(n16075), .B(n16074), .CI(n16073), .CO(n16086), .S(n16785)
         );
  ADDFHX1 U7341 ( .A(n9305), .B(n9304), .CI(n9303), .CO(n9314), .S(n9391) );
  INVX1 U7342 ( .A(n23207), .Y(n19354) );
  NAND2XL U7343 ( .A(n18590), .B(n18589), .Y(n6092) );
  ADDFHX1 U7344 ( .A(n12196), .B(n12195), .CI(n12194), .CO(n12410), .S(n12409)
         );
  NAND2X1 U7345 ( .A(n7388), .B(n7836), .Y(n7403) );
  OAI2BB1XL U7346 ( .A0N(n11890), .A1N(n4989), .B0(n4987), .Y(n11910) );
  NAND2XL U7347 ( .A(n17704), .B(n17703), .Y(n4336) );
  INVX1 U7348 ( .A(n21491), .Y(n21488) );
  ADDFHX1 U7349 ( .A(n17761), .B(n17760), .CI(n17759), .CO(n17797), .S(n17801)
         );
  OR2X2 U7350 ( .A(n24043), .B(n13003), .Y(n11604) );
  NAND2XL U7351 ( .A(n4934), .B(n3452), .Y(n4670) );
  NAND2X1 U7352 ( .A(n7674), .B(n7673), .Y(n7745) );
  NAND2X1 U7353 ( .A(n7675), .B(n7676), .Y(n7749) );
  ADDFHX1 U7354 ( .A(n12060), .B(n12059), .CI(n12058), .CO(n12440), .S(n12061)
         );
  INVXL U7355 ( .A(n12668), .Y(n5040) );
  ADDFHX1 U7356 ( .A(n7242), .B(n7241), .CI(n7240), .CO(n7121), .S(n7251) );
  XNOR2X1 U7357 ( .A(n10661), .B(M2_mult_x_15_n1668), .Y(n10662) );
  ADDFHX1 U7358 ( .A(n17064), .B(n17063), .CI(n17062), .CO(n17065), .S(n17051)
         );
  INVX1 U7359 ( .A(n16045), .Y(n4153) );
  XOR2X2 U7360 ( .A(n4956), .B(n11692), .Y(n3902) );
  OAI21X2 U7361 ( .A0(n15558), .A1(n14917), .B0(n14916), .Y(n24355) );
  INVXL U7362 ( .A(n18360), .Y(n4092) );
  NAND2XL U7363 ( .A(n17773), .B(n17774), .Y(n3752) );
  NAND2X1 U7364 ( .A(n4832), .B(n4831), .Y(n16171) );
  ADDFHX2 U7365 ( .A(n16802), .B(n16801), .CI(n16800), .CO(n16827), .S(n16831)
         );
  ADDFHX1 U7366 ( .A(n12402), .B(n12401), .CI(n12400), .CO(n12403), .S(n12380)
         );
  INVX1 U7367 ( .A(n20652), .Y(n4522) );
  OR2X2 U7368 ( .A(n20652), .B(n19025), .Y(n18766) );
  ADDFHX1 U7369 ( .A(n16260), .B(n16259), .CI(n16258), .CO(n16264), .S(n16244)
         );
  OAI22X1 U7370 ( .A0(n15559), .A1(n3101), .B0(n15558), .B1(n15557), .Y(n15570) );
  INVXL U7371 ( .A(n11719), .Y(n4428) );
  ADDFHX1 U7372 ( .A(n12369), .B(n12368), .CI(n12367), .CO(n12401), .S(n12370)
         );
  NAND2XL U7373 ( .A(n3041), .B(n19330), .Y(n19331) );
  OAI2BB1XL U7374 ( .A0N(n17939), .A1N(n4391), .B0(n4390), .Y(n17952) );
  NAND2BXL U7375 ( .AN(n13225), .B(n13173), .Y(n5165) );
  NAND2XL U7376 ( .A(n6769), .B(n6770), .Y(n3497) );
  NAND2X1 U7377 ( .A(n19564), .B(n19329), .Y(n19302) );
  NAND2X1 U7378 ( .A(n3041), .B(n19337), .Y(n19298) );
  OAI2BB1XL U7379 ( .A0N(n14250), .A1N(n14249), .B0(n14228), .Y(n14262) );
  NOR2X1 U7380 ( .A(n10676), .B(n10672), .Y(n9159) );
  NAND2X1 U7381 ( .A(n19566), .B(n19325), .Y(n19303) );
  NAND2XL U7382 ( .A(n18364), .B(n18363), .Y(n4193) );
  ADDFHX1 U7383 ( .A(n18285), .B(n18284), .CI(n18283), .CO(n18292), .S(n18291)
         );
  OAI21XL U7384 ( .A0(n17773), .A1(n17774), .B0(n17772), .Y(n3753) );
  XOR2X1 U7385 ( .A(n3381), .B(n5982), .Y(n12139) );
  ADDFHX1 U7386 ( .A(n7080), .B(n7079), .CI(n7078), .CO(n7242), .S(n7130) );
  INVXL U7387 ( .A(n14249), .Y(n3452) );
  ADDFHX1 U7388 ( .A(n12161), .B(n12160), .CI(n12159), .CO(n12156), .S(n12217)
         );
  OR2XL U7389 ( .A(n16656), .B(n16655), .Y(n16654) );
  INVX1 U7390 ( .A(n17594), .Y(n3098) );
  ADDFHX1 U7391 ( .A(n6999), .B(n6998), .CI(n6997), .CO(n7243), .S(n7002) );
  ADDFHX2 U7392 ( .A(n12116), .B(n12115), .CI(n12114), .CO(n12093), .S(n12137)
         );
  ADDFHX1 U7393 ( .A(n16741), .B(n16740), .CI(n16739), .CO(n16746), .S(n16748)
         );
  OAI21XL U7394 ( .A0(n5907), .A1(n5909), .B0(n5905), .Y(n17614) );
  ADDFHX2 U7395 ( .A(n18056), .B(n18055), .CI(n18054), .CO(n18097), .S(n18099)
         );
  ADDFHX1 U7396 ( .A(n18340), .B(n18339), .CI(n18338), .CO(n18355), .S(n18373)
         );
  NAND2XL U7397 ( .A(n3175), .B(n4074), .Y(n5413) );
  OAI21XL U7398 ( .A0(n11754), .A1(n11755), .B0(n11753), .Y(n3448) );
  INVXL U7399 ( .A(n10403), .Y(n4568) );
  NAND2XL U7400 ( .A(n15190), .B(n14943), .Y(n14944) );
  NAND2XL U7401 ( .A(n11694), .B(n11693), .Y(n4957) );
  AND2X2 U7402 ( .A(n17153), .B(n17152), .Y(n4702) );
  OAI21XL U7403 ( .A0(n7838), .A1(n7837), .B0(n7836), .Y(n23199) );
  NOR2X1 U7404 ( .A(n18759), .B(n19028), .Y(n19025) );
  NOR2X1 U7405 ( .A(n7698), .B(n7697), .Y(n7721) );
  NAND2X1 U7406 ( .A(n23406), .B(n21446), .Y(n21479) );
  ADDFHX1 U7407 ( .A(n11758), .B(n11757), .CI(n11756), .CO(n11868), .S(n11784)
         );
  OAI21X1 U7408 ( .A0(n16960), .A1(n5692), .B0(n5691), .Y(n16895) );
  NAND2XL U7409 ( .A(n5724), .B(n3176), .Y(n5723) );
  AND2X2 U7410 ( .A(n10660), .B(n10659), .Y(n10661) );
  XNOR3X2 U7411 ( .A(n6402), .B(n6401), .C(n3517), .Y(n6441) );
  NAND2X1 U7412 ( .A(n15190), .B(n14942), .Y(n14918) );
  NAND2X1 U7413 ( .A(n5824), .B(n3022), .Y(n17104) );
  ADDFHX1 U7414 ( .A(n7601), .B(n7600), .CI(n7599), .CO(n7603), .S(n7605) );
  ADDFHX1 U7415 ( .A(n12704), .B(n12703), .CI(n12702), .CO(n12705), .S(n12691)
         );
  NAND2XL U7416 ( .A(n3416), .B(n5782), .Y(n5779) );
  NAND2BXL U7417 ( .AN(n11891), .B(n4990), .Y(n4989) );
  INVX1 U7418 ( .A(n23122), .Y(n21446) );
  NOR2X1 U7419 ( .A(n10660), .B(M2_mult_x_15_n1668), .Y(n10570) );
  INVXL U7420 ( .A(n12707), .Y(n6000) );
  ADDFHX1 U7421 ( .A(n12393), .B(n12392), .CI(n12391), .CO(n12398), .S(n12400)
         );
  ADDFHX1 U7422 ( .A(n17911), .B(n17910), .CI(n17909), .CO(n17921), .S(n17918)
         );
  NAND3X1 U7423 ( .A(n23398), .B(n23420), .C(n23230), .Y(n21403) );
  INVX4 U7424 ( .A(n3041), .Y(n3100) );
  NAND4X1 U7425 ( .A(n23402), .B(n23394), .C(n23413), .D(n23406), .Y(n21404)
         );
  XOR2X1 U7426 ( .A(n17179), .B(n17400), .Y(n17186) );
  NOR2X1 U7427 ( .A(n9121), .B(n9120), .Y(n10672) );
  NAND2XL U7428 ( .A(n17092), .B(n17099), .Y(n5824) );
  ADDFHX1 U7429 ( .A(n6373), .B(n6372), .CI(n6371), .CO(n6386), .S(n6415) );
  NAND2X1 U7430 ( .A(n18711), .B(n18710), .Y(n19016) );
  OAI21XL U7431 ( .A0(n3929), .A1(n11833), .B0(n11832), .Y(n3926) );
  NAND2X1 U7432 ( .A(n18760), .B(n19029), .Y(n18759) );
  ADDFHX1 U7433 ( .A(n11956), .B(n11955), .CI(n11954), .CO(n11990), .S(n11959)
         );
  NAND2X1 U7434 ( .A(n18713), .B(n18712), .Y(n18996) );
  ADDFHX1 U7435 ( .A(n11945), .B(n11944), .CI(n11943), .CO(n11975), .S(n11960)
         );
  OR2XL U7436 ( .A(n12288), .B(n12287), .Y(n12286) );
  NAND2BXL U7437 ( .AN(n16287), .B(n3179), .Y(n5328) );
  OR2XL U7438 ( .A(n6586), .B(n6585), .Y(n6584) );
  INVX2 U7439 ( .A(n5414), .Y(n3175) );
  XOR2X1 U7440 ( .A(n3177), .B(n9904), .Y(n4303) );
  NAND2XL U7441 ( .A(n5982), .B(n3846), .Y(n5981) );
  BUFX2 U7442 ( .A(n16100), .Y(n4780) );
  NAND2X1 U7443 ( .A(n12998), .B(n12997), .Y(n12999) );
  XNOR2X1 U7444 ( .A(n9904), .B(n10386), .Y(n9706) );
  INVXL U7445 ( .A(n5546), .Y(n5545) );
  NAND2X1 U7446 ( .A(n7802), .B(n7801), .Y(n7816) );
  OAI2BB1XL U7447 ( .A0N(n4436), .A1N(n12541), .B0(n4435), .Y(n12549) );
  NOR2XL U7448 ( .A(n17720), .B(n3765), .Y(n3764) );
  ADDFHX1 U7449 ( .A(n11898), .B(n11897), .CI(n11896), .CO(n11931), .S(n11867)
         );
  XOR2X1 U7450 ( .A(n11754), .B(n11753), .Y(n3352) );
  ADDFHX1 U7451 ( .A(n17946), .B(n17945), .CI(n17944), .CO(n17961), .S(n17990)
         );
  NAND2XL U7452 ( .A(n3179), .B(n3952), .Y(n5946) );
  INVX1 U7453 ( .A(n10659), .Y(n10658) );
  NOR2XL U7454 ( .A(n9723), .B(n9694), .Y(n5748) );
  XOR2X1 U7455 ( .A(n10338), .B(n10341), .Y(n9252) );
  INVXL U7456 ( .A(n3440), .Y(n3439) );
  OR2XL U7457 ( .A(n18172), .B(n18171), .Y(n18170) );
  OR2XL U7458 ( .A(n12698), .B(n5996), .Y(n5994) );
  NAND3X1 U7459 ( .A(n9148), .B(n9147), .C(n14436), .Y(n10685) );
  NAND4X1 U7460 ( .A(n9131), .B(n9130), .C(n9129), .D(n25213), .Y(n10678) );
  ADDFHX1 U7461 ( .A(n18065), .B(n18064), .CI(n18063), .CO(n18058), .S(n18093)
         );
  XOR2X1 U7462 ( .A(M2_a_16_), .B(M2_a_17_), .Y(n5238) );
  NAND2XL U7463 ( .A(n6975), .B(n3561), .Y(n3560) );
  CLKINVX3 U7464 ( .A(n16962), .Y(n3179) );
  OAI2BB1XL U7465 ( .A0N(n16960), .A1N(n16962), .B0(n3211), .Y(n17041) );
  XOR2X1 U7466 ( .A(n6974), .B(n3563), .Y(n6960) );
  ADDFHX1 U7467 ( .A(n6987), .B(n6986), .CI(n6985), .CO(n7126), .S(n6983) );
  INVXL U7468 ( .A(n11833), .Y(n3927) );
  ADDFHX1 U7469 ( .A(n7303), .B(n7302), .CI(n7301), .CO(n7456), .S(n7274) );
  CLKINVX3 U7470 ( .A(n9843), .Y(n3282) );
  NAND2BXL U7471 ( .AN(n15965), .B(n3179), .Y(n3618) );
  AND2X2 U7472 ( .A(n17412), .B(n19042), .Y(n21170) );
  OAI22X1 U7473 ( .A0(n4039), .A1(n12119), .B0(n12618), .B1(n3875), .Y(n12076)
         );
  OR2XL U7474 ( .A(n16634), .B(n16633), .Y(n16632) );
  NAND2XL U7475 ( .A(n3874), .B(n3873), .Y(n3872) );
  ADDFHX1 U7476 ( .A(n6852), .B(n6853), .CI(n6854), .CO(n6884), .S(n6889) );
  ADDFHX1 U7477 ( .A(n6392), .B(n6391), .CI(n6390), .CO(n6384), .S(n6420) );
  ADDFHX1 U7478 ( .A(n12155), .B(n12154), .CI(n12153), .CO(n12161), .S(n12178)
         );
  AND2X1 U7479 ( .A(M4_U4_U1_enc_tree_3__3__16_), .B(
        M4_U4_U1_enc_tree_3__3__24_), .Y(n18810) );
  NOR2XL U7480 ( .A(n9901), .B(M2_b_2_), .Y(M2_U4_U1_enc_tree_1__1__28_) );
  NOR2XL U7481 ( .A(n9901), .B(n3182), .Y(M2_U4_U1_or2_tree_0__1__28_) );
  NAND2XL U7482 ( .A(n16974), .B(n4099), .Y(n4095) );
  NOR2XL U7483 ( .A(n11812), .B(n12759), .Y(n3656) );
  OR2X2 U7484 ( .A(n7832), .B(n7831), .Y(n7834) );
  OAI22X1 U7485 ( .A0(n21998), .A1(n3042), .B0(n3020), .B1(n21351), .Y(n22009)
         );
  ADDFHX1 U7486 ( .A(n16286), .B(n16285), .CI(n16284), .CO(n16326), .S(n16290)
         );
  XOR2X1 U7487 ( .A(n7391), .B(n7849), .Y(n7405) );
  NAND2XL U7488 ( .A(n5674), .B(n5642), .Y(n5641) );
  OAI22X1 U7489 ( .A0(n12357), .A1(n11671), .B0(n12284), .B1(n11652), .Y(
        n11684) );
  OAI2BB1X1 U7490 ( .A0N(n3451), .A1N(n3188), .B0(n5109), .Y(n7626) );
  NAND4X1 U7491 ( .A(n14456), .B(n14440), .C(n14439), .D(n14438), .Y(n14709)
         );
  NAND4X1 U7492 ( .A(n14456), .B(n14436), .C(n14435), .D(n14434), .Y(n14710)
         );
  INVX8 U7493 ( .A(n15008), .Y(n3101) );
  INVX4 U7494 ( .A(n19290), .Y(n19297) );
  OAI22XL U7495 ( .A0(n11629), .A1(n12715), .B0(n12525), .B1(n3350), .Y(n11630) );
  NAND2X1 U7496 ( .A(n18762), .B(n19032), .Y(n18761) );
  NAND2X1 U7497 ( .A(n3020), .B(n21435), .Y(n21436) );
  NAND2XL U7498 ( .A(n5898), .B(n3187), .Y(n5897) );
  XNOR2X1 U7499 ( .A(n12996), .B(n3202), .Y(n12997) );
  NAND3X1 U7500 ( .A(n9166), .B(n9165), .C(n14444), .Y(n10694) );
  NAND2X1 U7501 ( .A(n3020), .B(n21431), .Y(n21432) );
  NAND2BXL U7502 ( .AN(n16540), .B(n5847), .Y(n5842) );
  NAND3X1 U7503 ( .A(n9155), .B(n9154), .C(n14455), .Y(n10692) );
  NAND3X1 U7504 ( .A(n9151), .B(n9150), .C(n14440), .Y(n10687) );
  NAND2BXL U7505 ( .AN(n12095), .B(n5941), .Y(n4985) );
  OAI22X1 U7506 ( .A0(n12028), .A1(n12717), .B0(n12718), .B1(n3754), .Y(n12075) );
  OAI21XL U7507 ( .A0(n5460), .A1(n18107), .B0(n5459), .Y(n18017) );
  OAI22X1 U7508 ( .A0(n12715), .A1(n11814), .B0(n12525), .B1(n11744), .Y(n4926) );
  XNOR2X1 U7509 ( .A(n6975), .B(n3564), .Y(n3563) );
  OAI21XL U7510 ( .A0(n12152), .A1(n4008), .B0(n4007), .Y(n12146) );
  INVXL U7511 ( .A(n17939), .Y(n4031) );
  ADDFHX1 U7512 ( .A(n6743), .B(n6742), .CI(n6741), .CO(n6852), .S(n6763) );
  NAND2X1 U7513 ( .A(n21519), .B(n21426), .Y(n21427) );
  OAI21XL U7514 ( .A0(n12701), .A1(n3198), .B0(n3969), .Y(n3967) );
  NAND3X1 U7515 ( .A(n9158), .B(n9157), .C(n14448), .Y(n10695) );
  OAI22XL U7516 ( .A0(n12715), .A1(n6115), .B0(n12525), .B1(n11814), .Y(n11855) );
  INVXL U7517 ( .A(n12718), .Y(n5415) );
  OAI22XL U7518 ( .A0(n12099), .A1(n12598), .B0(n12065), .B1(n12342), .Y(n5980) );
  OAI2BB1XL U7519 ( .A0N(n12342), .A1N(n12598), .B0(n3204), .Y(n12631) );
  NAND2BXL U7520 ( .AN(n12125), .B(n3186), .Y(n6007) );
  OR2X4 U7521 ( .A(n14907), .B(n14906), .Y(n4467) );
  OAI22X1 U7522 ( .A0(n17148), .A1(n12701), .B0(n3194), .B1(n3198), .Y(n16908)
         );
  NAND2XL U7523 ( .A(n4165), .B(n4164), .Y(n4163) );
  NOR2X1 U7524 ( .A(n12535), .B(n3202), .Y(n12802) );
  NAND2BXL U7525 ( .AN(n7052), .B(n3188), .Y(n5120) );
  NAND2BXL U7526 ( .AN(n6977), .B(n3188), .Y(n5114) );
  NAND2BXL U7527 ( .AN(n7184), .B(n3188), .Y(n5117) );
  INVXL U7528 ( .A(n16942), .Y(n5732) );
  NAND2X1 U7529 ( .A(n14445), .B(n14697), .Y(n14441) );
  INVXL U7530 ( .A(n18107), .Y(n5458) );
  AOI21X1 U7531 ( .A0(n8157), .A1(n8156), .B0(n8155), .Y(n8158) );
  INVXL U7532 ( .A(n10159), .Y(n6065) );
  NAND2BXL U7533 ( .AN(n6345), .B(n3188), .Y(n5123) );
  NAND2X1 U7534 ( .A(n9059), .B(n11546), .Y(n9341) );
  INVXL U7535 ( .A(n12618), .Y(n4968) );
  NOR2X1 U7536 ( .A(n17148), .B(n3202), .Y(n17105) );
  XNOR2X1 U7537 ( .A(n17149), .B(n3202), .Y(n17150) );
  NAND4X1 U7538 ( .A(n13022), .B(n13021), .C(n13020), .D(n13019), .Y(n19042)
         );
  XNOR2X1 U7539 ( .A(n14358), .B(n14357), .Y(n14359) );
  OAI22XL U7540 ( .A0(n17941), .A1(n18239), .B0(n18141), .B1(n5815), .Y(n17939) );
  ADDFHX1 U7541 ( .A(n12271), .B(n11697), .CI(n11696), .CO(n11776), .S(n11699)
         );
  NAND2BXL U7542 ( .AN(n11637), .B(n3736), .Y(n3735) );
  NAND2XL U7543 ( .A(n4188), .B(n3192), .Y(n4186) );
  OAI21XL U7544 ( .A0(n7955), .A1(n7954), .B0(n7953), .Y(n8026) );
  NOR2X1 U7545 ( .A(n8002), .B(n8022), .Y(n8025) );
  NAND2BXL U7546 ( .AN(n17742), .B(n3193), .Y(n5928) );
  XOR2X1 U7547 ( .A(n18604), .B(n3043), .Y(n4249) );
  AND2X2 U7548 ( .A(n18721), .B(n17512), .Y(n18722) );
  NAND2BXL U7549 ( .AN(n18635), .B(n3193), .Y(n4199) );
  OR2XL U7550 ( .A(n3196), .B(n3048), .Y(n5052) );
  NAND2XL U7551 ( .A(n3196), .B(n3048), .Y(n5051) );
  INVX4 U7552 ( .A(n5676), .Y(n17099) );
  OAI22X1 U7553 ( .A0(n7149), .A1(n3046), .B0(n4592), .B1(n3542), .Y(n7160) );
  BUFX3 U7554 ( .A(M1_a_20_), .Y(n14307) );
  NOR2X1 U7555 ( .A(n2993), .B(n14357), .Y(n14305) );
  INVX1 U7556 ( .A(n14357), .Y(n14354) );
  BUFX3 U7557 ( .A(n12284), .Y(n3183) );
  NAND2X1 U7558 ( .A(n11536), .B(sigma10[9]), .Y(n3284) );
  NAND2X1 U7559 ( .A(n17183), .B(n17406), .Y(n17182) );
  NOR2X1 U7560 ( .A(n7829), .B(n25872), .Y(n7799) );
  INVX1 U7561 ( .A(n24359), .Y(n25222) );
  NAND2X1 U7562 ( .A(n19242), .B(n19285), .Y(n19288) );
  NAND2X1 U7563 ( .A(n11596), .B(n13013), .Y(n11592) );
  NOR2X1 U7564 ( .A(n8075), .B(n8133), .Y(n8113) );
  NAND2X1 U7565 ( .A(n18764), .B(n19035), .Y(n18763) );
  NAND2X1 U7566 ( .A(n7397), .B(n7841), .Y(n7395) );
  XOR2X1 U7567 ( .A(n18673), .B(n3205), .Y(n4169) );
  NAND2X1 U7568 ( .A(n11536), .B(learning_rate[5]), .Y(n3330) );
  INVXL U7569 ( .A(n16959), .Y(n3952) );
  ADDFHX1 U7570 ( .A(n7098), .B(n7097), .CI(n7096), .CO(n7137), .S(n7107) );
  AOI22XL U7571 ( .A0(n25754), .A1(sigma11[19]), .B0(sigma12[19]), .B1(n3024), 
        .Y(n20934) );
  OAI22X1 U7572 ( .A0(n12339), .A1(n12340), .B0(n12338), .B1(n4238), .Y(n12348) );
  BUFX3 U7573 ( .A(M1_a_0_), .Y(n13049) );
  INVXL U7574 ( .A(n18504), .Y(n3104) );
  NOR2XL U7575 ( .A(n18006), .B(n3206), .Y(M4_U3_U1_or2_tree_0__1__28_) );
  OAI211X1 U7576 ( .A0(n25898), .A1(n9087), .B0(n9057), .C0(n9056), .Y(n9058)
         );
  NOR2X1 U7577 ( .A(n19026), .B(n19027), .Y(n18764) );
  NAND2X1 U7578 ( .A(n8049), .B(n8122), .Y(n8075) );
  OAI21X2 U7579 ( .A0(n21392), .A1(n21391), .B0(n21390), .Y(n21393) );
  XOR2X1 U7580 ( .A(n12701), .B(n3198), .Y(n3968) );
  NAND2X1 U7581 ( .A(n8074), .B(n8131), .Y(n8133) );
  INVXL U7582 ( .A(n12616), .Y(n5941) );
  XOR2X1 U7583 ( .A(M5_a_6_), .B(n4785), .Y(n15948) );
  NOR2XL U7584 ( .A(n9087), .B(n25906), .Y(n5346) );
  XOR2X1 U7585 ( .A(n3048), .B(n6014), .Y(n17045) );
  BUFX3 U7586 ( .A(M1_a_3_), .Y(n13863) );
  NOR2XL U7587 ( .A(n3203), .B(n15968), .Y(M5_U3_U1_or2_tree_0__1__20_) );
  NOR2X1 U7588 ( .A(n17397), .B(n17398), .Y(n17183) );
  NOR2XL U7589 ( .A(n3200), .B(n5677), .Y(M5_U3_U1_enc_tree_1__1__12_) );
  XOR2X2 U7590 ( .A(n4795), .B(n3022), .Y(n15951) );
  NOR2X1 U7591 ( .A(n19172), .B(n19192), .Y(n19195) );
  INVXL U7592 ( .A(n7287), .Y(n3578) );
  XNOR2X1 U7593 ( .A(n3202), .B(M4_U3_U1_or2_inv_0__30_), .Y(n6035) );
  INVXL U7594 ( .A(n3197), .Y(n6146) );
  OAI21XL U7595 ( .A0(n14792), .A1(n14791), .B0(n14790), .Y(n14815) );
  NOR2X1 U7596 ( .A(n13004), .B(n13005), .Y(n11596) );
  NAND2X1 U7597 ( .A(n8001), .B(n8020), .Y(n8022) );
  NAND2X1 U7598 ( .A(n19171), .B(n19190), .Y(n19192) );
  AOI222XL U7599 ( .A0(n22953), .A1(n11071), .B0(n22897), .B1(n3218), .C0(
        n22952), .C1(n9109), .Y(n22620) );
  XOR2XL U7600 ( .A(n3211), .B(n6162), .Y(n15965) );
  XOR2X1 U7601 ( .A(n7286), .B(n3584), .Y(n7065) );
  AOI222XL U7602 ( .A0(n22953), .A1(n9109), .B0(n10797), .B1(n11074), .C0(
        n22952), .C1(n3219), .Y(n22687) );
  AOI222XL U7603 ( .A0(n23023), .A1(n9109), .B0(n22887), .B1(n11074), .C0(
        n23021), .C1(n3219), .Y(n22639) );
  AOI222XL U7604 ( .A0(n23023), .A1(n11062), .B0(n22887), .B1(n3217), .C0(
        n23021), .C1(n26493), .Y(n22956) );
  BUFX2 U7605 ( .A(n12560), .Y(n12518) );
  AOI21X1 U7606 ( .A0(n21389), .A1(n21388), .B0(n21387), .Y(n21390) );
  INVXL U7607 ( .A(n2978), .Y(n3207) );
  NAND2X1 U7608 ( .A(n19207), .B(n19251), .Y(n19220) );
  AOI222XL U7609 ( .A0(n23023), .A1(n11063), .B0(n22887), .B1(n23109), .C0(
        n23021), .C1(n11062), .Y(n22863) );
  INVX2 U7610 ( .A(M3_mult_x_15_b_1_), .Y(n11658) );
  NOR2XL U7611 ( .A(M4_a_17_), .B(n3757), .Y(M4_U3_U1_enc_tree_1__1__14_) );
  XOR2X1 U7612 ( .A(n5087), .B(n17038), .Y(n3395) );
  CLKBUFX8 U7613 ( .A(n25786), .Y(n25754) );
  OAI21XL U7614 ( .A0(n8005), .A1(n8004), .B0(n8003), .Y(n8010) );
  NOR2X1 U7615 ( .A(n8008), .B(n7977), .Y(n8011) );
  INVX1 U7616 ( .A(n3198), .Y(n3106) );
  CLKINVX3 U7617 ( .A(n12701), .Y(n3107) );
  OAI21X2 U7618 ( .A0(n26277), .A1(n15942), .B0(n3803), .Y(n4785) );
  NAND3X1 U7619 ( .A(n18752), .B(n18751), .C(n18750), .Y(n19032) );
  AND2XL U7620 ( .A(n25815), .B(y11[10]), .Y(n3820) );
  NOR2X1 U7621 ( .A(n8086), .B(n8138), .Y(n8098) );
  NAND3X1 U7622 ( .A(n17165), .B(n17164), .C(n17163), .Y(n17406) );
  AOI22XL U7623 ( .A0(n22486), .A1(sigma12[20]), .B0(n25750), .B1(sigma11[20]), 
        .Y(n24245) );
  NOR2X1 U7624 ( .A(n8060), .B(n8125), .Y(n8074) );
  NOR2X1 U7625 ( .A(n8037), .B(n8116), .Y(n8049) );
  NOR2XL U7626 ( .A(n3211), .B(n5646), .Y(M5_U3_U1_enc_tree_1__1__16_) );
  INVX8 U7627 ( .A(n6162), .Y(M3_mult_x_15_b_9_) );
  OR2XL U7628 ( .A(M4_a_19_), .B(M4_a_17_), .Y(M4_U3_U1_or2_tree_0__1__12_) );
  XNOR2X1 U7629 ( .A(n7621), .B(n3209), .Y(n3603) );
  NAND3X1 U7630 ( .A(n18746), .B(n18745), .C(n18744), .Y(n19035) );
  AOI222XL U7631 ( .A0(n22988), .A1(n11073), .B0(n22980), .B1(n11063), .C0(
        n22976), .C1(n23109), .Y(n22653) );
  AOI222XL U7632 ( .A0(n22932), .A1(n11071), .B0(n22904), .B1(n3218), .C0(
        n22931), .C1(n9109), .Y(n22625) );
  AOI222XL U7633 ( .A0(n22892), .A1(n23109), .B0(n22708), .B1(n11062), .C0(
        n22891), .C1(n3217), .Y(n22633) );
  AOI222XL U7634 ( .A0(n22988), .A1(n26493), .B0(n22980), .B1(n11059), .C0(
        n22976), .C1(n11058), .Y(n22855) );
  AOI222XL U7635 ( .A0(n22892), .A1(n11063), .B0(n22708), .B1(n23109), .C0(
        n22891), .C1(n11062), .Y(n22597) );
  AOI222XL U7636 ( .A0(n22928), .A1(n9109), .B0(n22700), .B1(n11074), .C0(
        n22927), .C1(n3219), .Y(n22544) );
  AOI222XL U7637 ( .A0(n23152), .A1(n11063), .B0(n23093), .B1(n23109), .C0(
        n23150), .C1(n11062), .Y(n23106) );
  BUFX3 U7638 ( .A(n11494), .Y(M3_mult_x_15_b_15_) );
  AOI222XL U7639 ( .A0(n22892), .A1(n3219), .B0(n22708), .B1(n11073), .C0(
        n22891), .C1(n11063), .Y(n22560) );
  AOI222XL U7640 ( .A0(n23152), .A1(n23109), .B0(n23093), .B1(n11062), .C0(
        n23150), .C1(n3217), .Y(n23110) );
  NOR2X1 U7641 ( .A(n7375), .B(n7374), .Y(n7839) );
  AOI222XL U7642 ( .A0(n22892), .A1(n11074), .B0(n22708), .B1(n3219), .C0(
        n22891), .C1(n11073), .Y(n22513) );
  AOI222XL U7643 ( .A0(n22892), .A1(n11073), .B0(n22708), .B1(n11063), .C0(
        n22891), .C1(n23109), .Y(n22571) );
  AOI222XL U7644 ( .A0(n23003), .A1(n26493), .B0(n22969), .B1(n11059), .C0(
        n23001), .C1(n11058), .Y(n22962) );
  AOI222XL U7645 ( .A0(n22928), .A1(n3220), .B0(n22700), .B1(n22867), .C0(
        n22927), .C1(n10775), .Y(n22741) );
  NAND3X1 U7646 ( .A(n11563), .B(n11562), .C(n11561), .Y(n13013) );
  AOI222XL U7647 ( .A0(n22988), .A1(n11059), .B0(n22980), .B1(n11058), .C0(
        n22976), .C1(n23151), .Y(n22691) );
  AOI222XL U7648 ( .A0(n23003), .A1(n11062), .B0(n22969), .B1(n3217), .C0(
        n23001), .C1(n26493), .Y(n22865) );
  AOI222XL U7649 ( .A0(n22892), .A1(n11062), .B0(n22708), .B1(n3217), .C0(
        n22891), .C1(n26493), .Y(n22812) );
  AOI222XL U7650 ( .A0(n22892), .A1(n3217), .B0(n22708), .B1(n23022), .C0(
        n22891), .C1(n11059), .Y(n22667) );
  AOI222XL U7651 ( .A0(n23152), .A1(n3219), .B0(n23093), .B1(n11073), .C0(
        n23150), .C1(n11063), .Y(n23100) );
  XNOR2X2 U7652 ( .A(M0_a_8_), .B(n3213), .Y(n3579) );
  AOI222XL U7653 ( .A0(n22988), .A1(n11074), .B0(n22980), .B1(n3219), .C0(
        n22976), .C1(n11073), .Y(n22675) );
  AOI222XL U7654 ( .A0(n23152), .A1(n9109), .B0(n23093), .B1(n11074), .C0(
        n23150), .C1(n3219), .Y(n23097) );
  AOI222XL U7655 ( .A0(n22928), .A1(n23109), .B0(n22700), .B1(n11062), .C0(
        n22927), .C1(n3217), .Y(n22753) );
  AOI222XL U7656 ( .A0(n22988), .A1(n9109), .B0(n22980), .B1(n11074), .C0(
        n22976), .C1(n3219), .Y(n22749) );
  AOI222XL U7657 ( .A0(n22892), .A1(n9109), .B0(n22708), .B1(n11074), .C0(
        n22891), .C1(n3219), .Y(n22535) );
  AOI222XL U7658 ( .A0(n23003), .A1(n11063), .B0(n22969), .B1(n23109), .C0(
        n23001), .C1(n11062), .Y(n22836) );
  AOI222XL U7659 ( .A0(n22928), .A1(n3219), .B0(n22700), .B1(n11073), .C0(
        n22927), .C1(n11063), .Y(n22793) );
  AOI222XL U7660 ( .A0(n23023), .A1(n11071), .B0(n22887), .B1(n3218), .C0(
        n23021), .C1(n9109), .Y(n22613) );
  AOI222XL U7661 ( .A0(n23152), .A1(n11073), .B0(n23093), .B1(n11063), .C0(
        n23150), .C1(n23109), .Y(n23103) );
  AOI222XL U7662 ( .A0(n23152), .A1(n26493), .B0(n23093), .B1(n11059), .C0(
        n23150), .C1(n11058), .Y(n23144) );
  AOI222XL U7663 ( .A0(n23003), .A1(n9109), .B0(n22969), .B1(n11074), .C0(
        n23001), .C1(n3219), .Y(n22616) );
  AOI222XL U7664 ( .A0(n22928), .A1(n3217), .B0(n22700), .B1(n23022), .C0(
        n22927), .C1(n11059), .Y(n22908) );
  AOI222XL U7665 ( .A0(n22928), .A1(n11074), .B0(n22700), .B1(n3219), .C0(
        n22927), .C1(n11073), .Y(n22502) );
  NAND2X1 U7666 ( .A(n14827), .B(n14871), .Y(n14840) );
  CLKINVX3 U7667 ( .A(n23174), .Y(n3214) );
  NOR2X1 U7668 ( .A(n19178), .B(n19158), .Y(n19181) );
  NOR2X1 U7669 ( .A(n8793), .B(n8315), .Y(n8119) );
  NAND2XL U7670 ( .A(n14417), .B(y11[19]), .Y(n3558) );
  NOR2X1 U7671 ( .A(n14779), .B(n14786), .Y(n14789) );
  NOR2X1 U7672 ( .A(n8167), .B(n8180), .Y(n8141) );
  NOR2X1 U7673 ( .A(n19165), .B(n19184), .Y(n19171) );
  NOR2X1 U7674 ( .A(n8691), .B(n8243), .Y(n8017) );
  NAND2X1 U7675 ( .A(n14740), .B(n14801), .Y(n14751) );
  NAND2X1 U7676 ( .A(n19219), .B(n19261), .Y(n19263) );
  BUFX12 U7677 ( .A(n2978), .Y(n3110) );
  NAND2BX2 U7678 ( .AN(M5_a_0_), .B(n15970), .Y(n16686) );
  NOR2X1 U7679 ( .A(n19201), .B(n19245), .Y(n19207) );
  OAI21X2 U7680 ( .A0(n26242), .A1(n25767), .B0(n5046), .Y(n5045) );
  NOR2BX2 U7681 ( .AN(n4969), .B(n4432), .Y(n4979) );
  NOR2X1 U7682 ( .A(n14845), .B(n14887), .Y(n14851) );
  OR2X2 U7683 ( .A(n4946), .B(n4929), .Y(n4945) );
  NOR2X1 U7684 ( .A(n14745), .B(n14804), .Y(n14750) );
  NOR2X1 U7685 ( .A(n19820), .B(n19373), .Y(n19187) );
  NOR2X1 U7686 ( .A(n14798), .B(n14739), .Y(n14801) );
  AOI222XL U7687 ( .A0(n22928), .A1(n11071), .B0(n22700), .B1(n3218), .C0(
        n22927), .C1(n9109), .Y(n22520) );
  AOI222XL U7688 ( .A0(n23152), .A1(n11071), .B0(n23093), .B1(n3218), .C0(
        n23150), .C1(n9109), .Y(n23094) );
  AOI222XL U7689 ( .A0(n22892), .A1(n11071), .B0(n22708), .B1(n3218), .C0(
        n22891), .C1(n9109), .Y(n22537) );
  NOR2X1 U7690 ( .A(n19810), .B(n19366), .Y(n19184) );
  AOI222XL U7691 ( .A0(n23152), .A1(n3218), .B0(n23093), .B1(n23089), .C0(
        n23150), .C1(n11074), .Y(n23090) );
  INVX1 U7692 ( .A(n8357), .Y(n8401) );
  NAND2XL U7693 ( .A(n19583), .B(n19554), .Y(n19118) );
  NAND2BX4 U7694 ( .AN(n10785), .B(n10784), .Y(n22912) );
  INVX2 U7695 ( .A(n20860), .Y(n25737) );
  BUFX3 U7696 ( .A(M0_b_8_), .Y(n7475) );
  OR2XL U7697 ( .A(n10799), .B(n11207), .Y(n22896) );
  BUFX3 U7698 ( .A(M0_b_11_), .Y(n25879) );
  NAND2BX4 U7699 ( .AN(n11207), .B(n10799), .Y(n22834) );
  AOI222XL U7700 ( .A0(n22928), .A1(n3218), .B0(n22700), .B1(n23089), .C0(
        n22927), .C1(n11074), .Y(n22509) );
  AOI222XL U7701 ( .A0(n22988), .A1(n3218), .B0(n22980), .B1(n23089), .C0(
        n22976), .C1(n11074), .Y(n22745) );
  AOI222XL U7702 ( .A0(n22988), .A1(n11071), .B0(n22980), .B1(n3218), .C0(
        n22976), .C1(n9109), .Y(n22573) );
  NAND2BX4 U7703 ( .AN(n10760), .B(n10759), .Y(n23025) );
  BUFX3 U7704 ( .A(M0_b_6_), .Y(n25882) );
  NOR2BX4 U7705 ( .AN(n10760), .B(n10758), .Y(n22887) );
  AOI21X1 U7706 ( .A0(n4875), .A1(data[48]), .B0(n5420), .Y(n5419) );
  NOR2X1 U7707 ( .A(n14832), .B(n14874), .Y(n14839) );
  INVX1 U7708 ( .A(n8235), .Y(n8674) );
  INVX4 U7709 ( .A(n25813), .Y(n3111) );
  AND2XL U7710 ( .A(n5015), .B(data[124]), .Y(n17174) );
  INVX1 U7711 ( .A(n8316), .Y(n8793) );
  INVX1 U7712 ( .A(n8309), .Y(n8772) );
  NAND2X1 U7713 ( .A(n21349), .B(n21302), .Y(n21315) );
  NOR2X1 U7714 ( .A(n4531), .B(n4530), .Y(n4529) );
  INVX1 U7715 ( .A(n8307), .Y(n8712) );
  NOR2X1 U7716 ( .A(n19299), .B(n4803), .Y(n19230) );
  NOR2X1 U7717 ( .A(n14913), .B(n14926), .Y(n14890) );
  NOR2X1 U7718 ( .A(n19225), .B(n19268), .Y(n19231) );
  NAND2X2 U7719 ( .A(n11542), .B(n11541), .Y(M1_b_19_) );
  INVX1 U7720 ( .A(n8313), .Y(n8788) );
  NAND3X1 U7721 ( .A(n7377), .B(n7376), .C(n14410), .Y(n7841) );
  INVX1 U7722 ( .A(n8244), .Y(n8691) );
  INVX1 U7723 ( .A(n8261), .Y(n8659) );
  NAND2XL U7724 ( .A(n21231), .B(n21218), .Y(n21233) );
  AOI21XL U7725 ( .A0(n21231), .A1(n21230), .B0(n21229), .Y(n21232) );
  OAI21X2 U7726 ( .A0(n25767), .A1(n26257), .B0(n4895), .Y(n11480) );
  OAI2BB1X1 U7727 ( .A0N(y10[27]), .A1N(n3224), .B0(n7394), .Y(n7854) );
  OAI2BB1X1 U7728 ( .A0N(y10[23]), .A1N(n3224), .B0(n7401), .Y(n7858) );
  INVX1 U7729 ( .A(n8256), .Y(n8349) );
  NOR2X1 U7730 ( .A(n4539), .B(n4538), .Y(n4537) );
  OAI2BB1X1 U7731 ( .A0N(y10[28]), .A1N(n3224), .B0(n7392), .Y(n7855) );
  AND2X2 U7732 ( .A(n9066), .B(n3259), .Y(n3258) );
  NOR2X1 U7733 ( .A(n14821), .B(n14865), .Y(n14827) );
  CLKINVX3 U7734 ( .A(n25786), .Y(n25255) );
  CLKINVX3 U7735 ( .A(n3117), .Y(n4575) );
  NAND2BX4 U7736 ( .AN(n21082), .B(n21081), .Y(n23005) );
  INVX1 U7737 ( .A(n19487), .Y(n19532) );
  INVX1 U7738 ( .A(n15106), .Y(n15150) );
  NOR2BX4 U7739 ( .AN(n21082), .B(n21080), .Y(n22969) );
  NAND2XL U7740 ( .A(n5480), .B(sigma11[6]), .Y(n5892) );
  INVX1 U7741 ( .A(n19393), .Y(n19794) );
  INVX1 U7742 ( .A(n19386), .Y(n19479) );
  NOR2XL U7743 ( .A(n21223), .B(n21217), .Y(n21218) );
  NAND2BX4 U7744 ( .AN(n22563), .B(n22562), .Y(n22984) );
  NOR2BX4 U7745 ( .AN(n22563), .B(n21064), .Y(n22980) );
  INVXL U7746 ( .A(n19561), .Y(n19720) );
  INVX1 U7747 ( .A(n19371), .Y(n19815) );
  NOR2X1 U7748 ( .A(n14911), .B(n14930), .Y(n14856) );
  NOR2X1 U7749 ( .A(n15430), .B(n14982), .Y(n14804) );
  INVX1 U7750 ( .A(n19367), .Y(n19810) );
  NOR2X1 U7751 ( .A(n19922), .B(n19444), .Y(n19248) );
  INVX1 U7752 ( .A(n14955), .Y(n14915) );
  NOR2X1 U7753 ( .A(n15542), .B(n15065), .Y(n14868) );
  NOR2BX4 U7754 ( .AN(n22512), .B(n22493), .Y(n22708) );
  NAND2BX4 U7755 ( .AN(n22512), .B(n22511), .Y(n22894) );
  NOR2X1 U7756 ( .A(n15552), .B(n15049), .Y(n14874) );
  NOR2BX4 U7757 ( .AN(n21057), .B(n11090), .Y(n23093) );
  NOR2X1 U7758 ( .A(n15537), .B(n15062), .Y(n14826) );
  AOI22X1 U7759 ( .A0(n5480), .A1(sigma11[16]), .B0(in_valid_t), .B1(w2[48]), 
        .Y(n17475) );
  NOR2X1 U7760 ( .A(n15521), .B(n15058), .Y(n14865) );
  NAND2BX4 U7761 ( .AN(n21072), .B(n21071), .Y(n22909) );
  NOR2BX4 U7762 ( .AN(n21072), .B(n21070), .Y(n22700) );
  INVX1 U7763 ( .A(n19436), .Y(n19841) );
  INVXL U7764 ( .A(n19568), .Y(n19752) );
  INVX1 U7765 ( .A(n19365), .Y(n19802) );
  NOR2X1 U7766 ( .A(n19296), .B(n19310), .Y(n19271) );
  NOR2X1 U7767 ( .A(n21313), .B(n21354), .Y(n21314) );
  NOR2X1 U7768 ( .A(n21257), .B(n21277), .Y(n21258) );
  NAND4X1 U7769 ( .A(n8046), .B(n8045), .C(n8044), .D(n8043), .Y(n8313) );
  NAND4X1 U7770 ( .A(n8035), .B(n8034), .C(n8033), .D(n8032), .Y(n8309) );
  NAND4X1 U7771 ( .A(n7970), .B(n7969), .C(n7968), .D(n7967), .Y(n8264) );
  NAND4X1 U7772 ( .A(n7998), .B(n7997), .C(n7996), .D(n7995), .Y(n8241) );
  NAND4X1 U7773 ( .A(n8030), .B(n8029), .C(n8028), .D(n8027), .Y(n8307) );
  NAND2XL U7774 ( .A(n21166), .B(sigma12[8]), .Y(n5728) );
  INVX1 U7775 ( .A(n14998), .Y(n15097) );
  NOR2X1 U7776 ( .A(n21338), .B(n21517), .Y(n21341) );
  NAND2XL U7777 ( .A(n21350), .B(n21509), .Y(n21353) );
  NAND2XL U7778 ( .A(n21337), .B(n21514), .Y(n21340) );
  NOR2BXL U7779 ( .AN(n21166), .B(n6215), .Y(n4822) );
  NAND2X1 U7780 ( .A(n8104), .B(y20[29]), .Y(n8105) );
  NOR2XL U7781 ( .A(n21355), .B(n21421), .Y(n21307) );
  CLKINVX4 U7782 ( .A(n26494), .Y(n3220) );
  AOI22X1 U7783 ( .A0(n7389), .A1(target_temp[20]), .B0(in_valid_d), .B1(
        w1[20]), .Y(n6257) );
  INVX1 U7784 ( .A(n15059), .Y(n15521) );
  XNOR2X1 U7785 ( .A(n3058), .B(n22491), .Y(n22512) );
  AND2X2 U7786 ( .A(n21380), .B(n21417), .Y(n21381) );
  INVX1 U7787 ( .A(n14989), .Y(n15440) );
  NAND2XL U7788 ( .A(n7389), .B(y10[14]), .Y(n3477) );
  NAND2X1 U7789 ( .A(n5604), .B(w2[13]), .Y(n3478) );
  INVX1 U7790 ( .A(n15002), .Y(n15406) );
  INVX1 U7791 ( .A(n15063), .Y(n15537) );
  NAND2XL U7792 ( .A(n21265), .B(n21475), .Y(n21268) );
  INVX1 U7793 ( .A(n15057), .Y(n15461) );
  NAND2X1 U7794 ( .A(n21166), .B(sigma12[21]), .Y(n6017) );
  INVX2 U7795 ( .A(n11499), .Y(n3114) );
  XOR2X2 U7796 ( .A(n23202), .B(n23201), .Y(n19952) );
  NAND2XL U7797 ( .A(n21219), .B(n21604), .Y(n21222) );
  NOR2XL U7798 ( .A(n21278), .B(n21461), .Y(n21251) );
  INVX1 U7799 ( .A(n19442), .Y(n19917) );
  CLKBUFX3 U7800 ( .A(n11143), .Y(n11074) );
  NAND2XL U7801 ( .A(n21273), .B(n21457), .Y(n21276) );
  INVX1 U7802 ( .A(n11141), .Y(n26490) );
  NAND2X1 U7803 ( .A(n21166), .B(target_temp[10]), .Y(n6149) );
  CLKINVX3 U7804 ( .A(n22621), .Y(n3221) );
  NOR2XL U7805 ( .A(n21219), .B(n21604), .Y(n21217) );
  NOR2BX4 U7806 ( .AN(n10785), .B(n10783), .Y(n22904) );
  OAI21X1 U7807 ( .A0(n14833), .A1(n26515), .B0(n8091), .Y(n8180) );
  NAND2XL U7808 ( .A(n21366), .B(n21430), .Y(n21369) );
  INVX2 U7809 ( .A(n11133), .Y(n11395) );
  INVX1 U7810 ( .A(n14981), .Y(n15422) );
  INVXL U7811 ( .A(n21600), .Y(n21224) );
  NAND2XL U7812 ( .A(n3224), .B(y10[19]), .Y(n3585) );
  OAI21XL U7813 ( .A0(n3063), .A1(n25966), .B0(n4466), .Y(n14987) );
  INVXL U7814 ( .A(n21578), .Y(n21220) );
  OR2XL U7815 ( .A(n23884), .B(n26566), .Y(n4714) );
  BUFX2 U7816 ( .A(n11160), .Y(n10769) );
  BUFX2 U7817 ( .A(n11162), .Y(n10775) );
  BUFX2 U7818 ( .A(n11155), .Y(n10789) );
  OAI21X1 U7819 ( .A0(n3063), .A1(n19351), .B0(n19350), .Y(n23201) );
  XNOR2X1 U7820 ( .A(n23117), .B(n23115), .Y(n21527) );
  OR2XL U7821 ( .A(n23884), .B(n26559), .Y(n4713) );
  INVX1 U7822 ( .A(n23022), .Y(n26492) );
  INVX1 U7823 ( .A(n21977), .Y(n21338) );
  INVXL U7824 ( .A(n21844), .Y(n21261) );
  INVXL U7825 ( .A(n21809), .Y(n21201) );
  INVX8 U7826 ( .A(n21113), .Y(n3117) );
  NAND2X1 U7827 ( .A(n6217), .B(y10[30]), .Y(n7889) );
  INVX4 U7828 ( .A(n4710), .Y(n3118) );
  INVX8 U7829 ( .A(n9146), .Y(n3223) );
  AOI22X1 U7830 ( .A0(y12[23]), .A1(n19349), .B0(n3026), .B1(temp3[23]), .Y(
        n14835) );
  OR2XL U7831 ( .A(n21194), .B(n21620), .Y(n21184) );
  AOI22X1 U7832 ( .A0(y12[29]), .A1(n19349), .B0(n19216), .B1(temp3[29]), .Y(
        n14855) );
  AOI22X1 U7833 ( .A0(w2[94]), .A1(n19349), .B0(n3026), .B1(w1[126]), .Y(
        n14857) );
  INVX4 U7834 ( .A(n21112), .Y(n3226) );
  OAI21XL U7835 ( .A0(n26180), .A1(n21256), .B0(n21208), .Y(n21530) );
  CLKINVX8 U7836 ( .A(n3059), .Y(n3120) );
  AOI22X1 U7837 ( .A0(y10[23]), .A1(n19235), .B0(n3062), .B1(temp1[23]), .Y(
        n8065) );
  CLKINVX3 U7838 ( .A(n25693), .Y(n6161) );
  NAND2X1 U7839 ( .A(n11086), .B(n11085), .Y(n11210) );
  NAND2X1 U7840 ( .A(n21331), .B(temp0[31]), .Y(n21443) );
  INVX4 U7841 ( .A(n26595), .Y(n19349) );
  CLKINVX3 U7842 ( .A(n26595), .Y(n19235) );
  NAND2X1 U7843 ( .A(n21329), .B(temp0[24]), .Y(n21304) );
  NAND2XL U7844 ( .A(n21311), .B(w1[17]), .Y(n21297) );
  INVX4 U7845 ( .A(n21111), .Y(n19216) );
  NAND2XL U7846 ( .A(n21329), .B(w1[25]), .Y(n21321) );
  NAND2XL U7847 ( .A(n21331), .B(w1[10]), .Y(n21240) );
  NAND2XL U7848 ( .A(n21331), .B(w1[4]), .Y(n21173) );
  NAND2XL U7849 ( .A(n21311), .B(w1[5]), .Y(n21215) );
  NAND2X4 U7850 ( .A(n4584), .B(n4143), .Y(n9146) );
  NAND2XL U7851 ( .A(n21329), .B(w1[15]), .Y(n21249) );
  NAND2XL U7852 ( .A(n21333), .B(w1[16]), .Y(n21247) );
  CLKBUFX8 U7853 ( .A(n7881), .Y(n25693) );
  NAND2X1 U7854 ( .A(n11185), .B(n11184), .Y(n22990) );
  NAND2XL U7855 ( .A(n21311), .B(w1[20]), .Y(n21292) );
  NAND2XL U7856 ( .A(n21311), .B(w1[12]), .Y(n21235) );
  NAND2XL U7857 ( .A(n21329), .B(w1[27]), .Y(n21318) );
  NAND2XL U7858 ( .A(n21329), .B(w1[6]), .Y(n21213) );
  NAND2X1 U7859 ( .A(n21331), .B(temp0[30]), .Y(n21328) );
  NAND2X1 U7860 ( .A(n21329), .B(w1[29]), .Y(n21330) );
  NAND2XL U7861 ( .A(n21329), .B(w1[8]), .Y(n21208) );
  NAND2XL U7862 ( .A(n21329), .B(w1[7]), .Y(n21210) );
  NOR2X2 U7863 ( .A(n25542), .B(n21111), .Y(n21112) );
  NAND2X1 U7864 ( .A(n21331), .B(temp0[29]), .Y(n21332) );
  INVX8 U7865 ( .A(n25807), .Y(n3121) );
  INVX8 U7866 ( .A(n3228), .Y(n25567) );
  CLKINVX8 U7867 ( .A(n3228), .Y(n23088) );
  AND2X1 U7868 ( .A(n23973), .B(n26213), .Y(n5582) );
  OR2X4 U7869 ( .A(n7882), .B(n25886), .Y(n4637) );
  INVX4 U7870 ( .A(n4631), .Y(n21331) );
  INVX4 U7871 ( .A(n24632), .Y(n3122) );
  INVX1 U7872 ( .A(n25156), .Y(n4770) );
  MXI2XL U7873 ( .A(data[94]), .B(data[126]), .S0(n3229), .Y(n1708) );
  INVXL U7874 ( .A(n25145), .Y(n3259) );
  NAND2X1 U7875 ( .A(in_valid_d), .B(data_point[26]), .Y(n14410) );
  MXI2XL U7876 ( .A(data[88]), .B(data[120]), .S0(n3229), .Y(n1702) );
  MXI2XL U7877 ( .A(data[90]), .B(data[122]), .S0(n3229), .Y(n1704) );
  NAND2XL U7878 ( .A(in_valid_d), .B(w1[130]), .Y(n4550) );
  NAND2X1 U7879 ( .A(in_valid_t), .B(learning_rate[27]), .Y(n11585) );
  NAND2X1 U7880 ( .A(in_valid_t), .B(learning_rate[29]), .Y(n11577) );
  NAND2X1 U7881 ( .A(in_valid_t), .B(learning_rate[23]), .Y(n11600) );
  AND2X2 U7882 ( .A(in_valid_t), .B(w2[53]), .Y(n6094) );
  XNOR2X1 U7883 ( .A(cs[0]), .B(cs[1]), .Y(n7882) );
  NAND2X1 U7884 ( .A(in_valid_t), .B(learning_rate[5]), .Y(n6010) );
  NAND2XL U7885 ( .A(n4581), .B(data[115]), .Y(n3556) );
  NOR2X1 U7886 ( .A(n4585), .B(n6238), .Y(n25156) );
  INVX1 U7887 ( .A(data_point[18]), .Y(n6238) );
  INVX1 U7888 ( .A(data_point[5]), .Y(n6242) );
  INVX1 U7889 ( .A(data_point[20]), .Y(n6255) );
  INVX1 U7890 ( .A(data_point[10]), .Y(n6225) );
  INVX8 U7891 ( .A(n4586), .Y(n3123) );
  INVX1 U7892 ( .A(data_point[12]), .Y(n6250) );
  INVX1 U7893 ( .A(data_point[8]), .Y(n6263) );
  INVX1 U7894 ( .A(data_point[9]), .Y(n6227) );
  INVX8 U7895 ( .A(in_valid_t), .Y(n3398) );
  INVX1 U7896 ( .A(data_point[1]), .Y(n6277) );
  NAND3X1 U7897 ( .A(n24464), .B(n3315), .C(n3314), .Y(n24465) );
  INVX1 U7898 ( .A(n24652), .Y(n25495) );
  AOI21XL U7899 ( .A0(n23837), .A1(n25737), .B0(n4813), .Y(n2379) );
  AOI22X1 U7900 ( .A0(n24692), .A1(n24630), .B0(n24908), .B1(n24629), .Y(
        n24631) );
  OAI2BB1XL U7901 ( .A0N(n25741), .A1N(n25372), .B0(n5558), .Y(n5557) );
  OAI21XL U7902 ( .A0(n25535), .A1(n4571), .B0(n25534), .Y(n2040) );
  AOI22XL U7903 ( .A0(n24692), .A1(n24577), .B0(n24908), .B1(n24576), .Y(
        n24578) );
  AOI222XL U7904 ( .A0(n25735), .A1(n25737), .B0(n25743), .B1(y20[15]), .C0(
        n25734), .C1(n20890), .Y(n2375) );
  INVXL U7905 ( .A(n24374), .Y(n25262) );
  OAI21XL U7906 ( .A0(n25685), .A1(n3057), .B0(n25684), .Y(n25686) );
  INVX1 U7907 ( .A(n23577), .Y(n25520) );
  AOI222XL U7908 ( .A0(n25224), .A1(n25292), .B0(in_valid_w2), .B1(weight2[24]), .C0(w2[88]), .C1(n25822), .Y(n2224) );
  AOI22X1 U7909 ( .A0(n20385), .A1(n20864), .B0(n25300), .B1(n20863), .Y(
        n23577) );
  INVX1 U7910 ( .A(n25120), .Y(n25224) );
  AOI22X1 U7911 ( .A0(n20385), .A1(n23754), .B0(n25300), .B1(n23753), .Y(
        n23756) );
  NAND2X1 U7912 ( .A(n4450), .B(n4449), .Y(n24374) );
  NAND2X1 U7913 ( .A(n20234), .B(n20994), .Y(n24813) );
  AND2XL U7914 ( .A(n25284), .B(n25283), .Y(n25285) );
  AOI222X1 U7915 ( .A0(n24100), .A1(n24430), .B0(n24099), .B1(n24428), .C0(
        n24427), .C1(n24098), .Y(n25120) );
  AOI222X1 U7916 ( .A0(n24020), .A1(n24430), .B0(n24019), .B1(n24428), .C0(
        n24427), .C1(n24018), .Y(n25853) );
  AOI222X1 U7917 ( .A0(n24355), .A1(n24430), .B0(n24354), .B1(n24428), .C0(
        n24427), .C1(n24353), .Y(n24363) );
  AOI22XL U7918 ( .A0(n24427), .A1(n24058), .B0(n24430), .B1(n4787), .Y(n4449)
         );
  NAND2X1 U7919 ( .A(n24070), .B(n20169), .Y(n20172) );
  INVX1 U7920 ( .A(n24516), .Y(n24586) );
  INVXL U7921 ( .A(n23260), .Y(n2232) );
  NOR2X1 U7922 ( .A(n20233), .B(n24476), .Y(n20994) );
  NAND2X1 U7923 ( .A(n20516), .B(n20848), .Y(n20529) );
  NOR2X1 U7924 ( .A(n24646), .B(n20262), .Y(n24811) );
  AND2X2 U7925 ( .A(n23959), .B(n23961), .Y(n24427) );
  NAND2X1 U7926 ( .A(n15902), .B(n24516), .Y(n15935) );
  OR2X2 U7927 ( .A(n23961), .B(n23962), .Y(n4451) );
  NAND2X1 U7928 ( .A(n23959), .B(n15785), .Y(n15793) );
  NOR2X1 U7929 ( .A(n24658), .B(n15871), .Y(n24667) );
  INVXL U7930 ( .A(n24950), .Y(n24905) );
  INVX1 U7931 ( .A(n23312), .Y(n23359) );
  INVXL U7932 ( .A(n24808), .Y(n24728) );
  INVX1 U7933 ( .A(n23375), .Y(n23389) );
  INVX1 U7934 ( .A(n23271), .Y(n23364) );
  INVX1 U7935 ( .A(n23276), .Y(n23363) );
  INVX1 U7936 ( .A(n23381), .Y(n23390) );
  INVX1 U7937 ( .A(n23317), .Y(n23360) );
  INVX1 U7938 ( .A(n23291), .Y(n23365) );
  NOR2X1 U7939 ( .A(n15901), .B(n24482), .Y(n24516) );
  INVXL U7940 ( .A(n24663), .Y(n24660) );
  INVX1 U7941 ( .A(n23323), .Y(n23361) );
  AND2XL U7942 ( .A(n23798), .B(n20603), .Y(n20604) );
  INVX1 U7943 ( .A(n23336), .Y(n23366) );
  INVX1 U7944 ( .A(n23328), .Y(n23362) );
  INVX1 U7945 ( .A(n23388), .Y(n23391) );
  INVX1 U7946 ( .A(n23351), .Y(n23368) );
  INVX1 U7947 ( .A(n23247), .Y(n23249) );
  NAND2XL U7948 ( .A(n24686), .B(n24685), .Y(n24687) );
  INVX1 U7949 ( .A(n23342), .Y(n23367) );
  NAND2X1 U7950 ( .A(n20528), .B(n20884), .Y(n20838) );
  INVX1 U7951 ( .A(n23266), .Y(n23352) );
  INVX1 U7952 ( .A(n23306), .Y(n23358) );
  INVX1 U7953 ( .A(n23298), .Y(n23357) );
  INVX1 U7954 ( .A(n23243), .Y(n23248) );
  INVX1 U7955 ( .A(n4781), .Y(n4782) );
  INVX1 U7956 ( .A(n20884), .Y(n24562) );
  INVX1 U7957 ( .A(n23286), .Y(n23353) );
  INVX1 U7958 ( .A(n23283), .Y(n23354) );
  NOR2X1 U7959 ( .A(n15870), .B(n15869), .Y(n24663) );
  NAND2X2 U7960 ( .A(n4452), .B(n4617), .Y(n23963) );
  NOR2X1 U7961 ( .A(n24299), .B(n20128), .Y(n20134) );
  NOR2X1 U7962 ( .A(n20901), .B(n20515), .Y(n20848) );
  NOR2X1 U7963 ( .A(n20527), .B(n20909), .Y(n20884) );
  NOR2X1 U7964 ( .A(n20193), .B(n20192), .Y(n24725) );
  AOI222XL U7965 ( .A0(n23422), .A1(n23429), .B0(target_temp[26]), .B1(n23428), 
        .C0(in_valid_t), .C1(target[26]), .Y(n2258) );
  AOI222XL U7966 ( .A0(n23425), .A1(n23429), .B0(target_temp[23]), .B1(n23428), 
        .C0(in_valid_t), .C1(target[23]), .Y(n2255) );
  OR3X2 U7967 ( .A(n24019), .B(n24429), .C(n15750), .Y(n4617) );
  NOR2X1 U7968 ( .A(n15842), .B(n15841), .Y(n24622) );
  NOR2X1 U7969 ( .A(n15887), .B(n15886), .Y(n24670) );
  NOR2X1 U7970 ( .A(n24756), .B(n23200), .Y(n20154) );
  AOI222XL U7971 ( .A0(n23426), .A1(n23429), .B0(target_temp[29]), .B1(n23428), 
        .C0(in_valid_t), .C1(target[29]), .Y(n2261) );
  AOI222XL U7972 ( .A0(n23424), .A1(n23429), .B0(target_temp[28]), .B1(n23428), 
        .C0(in_valid_t), .C1(target[28]), .Y(n2260) );
  NOR2X1 U7973 ( .A(n15880), .B(n15879), .Y(n24703) );
  AOI222XL U7974 ( .A0(n23430), .A1(n23429), .B0(target_temp[25]), .B1(n23428), 
        .C0(in_valid_t), .C1(target[25]), .Y(n2257) );
  AOI222XL U7975 ( .A0(n23427), .A1(n23429), .B0(target_temp[24]), .B1(n23428), 
        .C0(in_valid_t), .C1(target[24]), .Y(n2256) );
  NOR2BX1 U7976 ( .AN(n20132), .B(n20131), .Y(n20133) );
  AOI222XL U7977 ( .A0(n23423), .A1(n25541), .B0(n4576), .B1(w1[286]), .C0(
        n23088), .C1(w1[318]), .Y(n2131) );
  AOI2BB1X1 U7978 ( .A0N(n20066), .A1N(n24848), .B0(n20253), .Y(n24630) );
  AOI222XL U7979 ( .A0(n23423), .A1(n23429), .B0(target_temp[30]), .B1(n23428), 
        .C0(in_valid_t), .C1(target[30]), .Y(n2262) );
  AOI2BB1X1 U7980 ( .A0N(n20066), .A1N(n24797), .B0(n20247), .Y(n24607) );
  NAND2XL U7981 ( .A(n20429), .B(n20428), .Y(n20430) );
  AOI2BB1X1 U7982 ( .A0N(n15688), .A1N(n24869), .B0(n15855), .Y(n24637) );
  OAI22XL U7983 ( .A0(n15891), .A1(n15688), .B0(n15890), .B1(n3077), .Y(n25280) );
  OAI21XL U7984 ( .A0(n23233), .A1(n23232), .B0(n23231), .Y(n23234) );
  AOI2BB1X1 U7985 ( .A0N(n15688), .A1N(n15909), .B0(n15850), .Y(n24618) );
  NOR2BX1 U7986 ( .AN(n15738), .B(n15737), .Y(n15751) );
  NAND2X1 U7987 ( .A(n20246), .B(n3075), .Y(n24804) );
  NAND2X1 U7988 ( .A(n20225), .B(n3075), .Y(n24756) );
  NAND2XL U7989 ( .A(n3077), .B(n15888), .Y(n25019) );
  NAND2X1 U7990 ( .A(n20216), .B(n3075), .Y(n24722) );
  NAND2X1 U7991 ( .A(n15919), .B(n3076), .Y(n15769) );
  NOR2X1 U7992 ( .A(n20230), .B(n20182), .Y(n20225) );
  NOR2XL U7993 ( .A(n15877), .B(n15808), .Y(n15900) );
  NOR2X1 U7994 ( .A(n20208), .B(n20207), .Y(n20232) );
  NOR2X1 U7995 ( .A(n20228), .B(n20182), .Y(n20216) );
  NOR3X1 U7996 ( .A(n24435), .B(n24391), .C(n20121), .Y(n20129) );
  AOI2BB1X1 U7997 ( .A0N(n20597), .A1N(n20572), .B0(n20514), .Y(n20877) );
  NOR2BXL U7998 ( .AN(n15739), .B(n24018), .Y(n15738) );
  OAI22XL U7999 ( .A0(n20590), .A1(n3073), .B0(n20589), .B1(n20588), .Y(n23805) );
  AOI2BB1X1 U8000 ( .A0N(n20522), .A1N(n20597), .B0(n20521), .Y(n20889) );
  OR2XL U8001 ( .A(n20427), .B(n20576), .Y(n20428) );
  NOR2X1 U8002 ( .A(n20480), .B(n20479), .Y(n24712) );
  NOR2X1 U8003 ( .A(n20466), .B(n8997), .Y(n9013) );
  AOI2BB1X1 U8004 ( .A0N(n20597), .A1N(n20537), .B0(n20503), .Y(n23583) );
  NOR2X1 U8005 ( .A(n15894), .B(n15688), .Y(n15919) );
  NAND3BX1 U8006 ( .AN(n9008), .B(n20431), .C(n9007), .Y(n9014) );
  NAND2X1 U8007 ( .A(n20520), .B(n20576), .Y(n20466) );
  NOR2X1 U8008 ( .A(n20498), .B(n20497), .Y(n20864) );
  XOR2X1 U8009 ( .A(n15742), .B(n15741), .Y(n24400) );
  AND2X2 U8010 ( .A(n23228), .B(n4768), .Y(n23418) );
  NOR2BXL U8011 ( .AN(n8991), .B(n23691), .Y(n8994) );
  NAND2X1 U8012 ( .A(n20395), .B(n20576), .Y(n20431) );
  NOR2XL U8013 ( .A(n20465), .B(n20464), .Y(n20467) );
  AND2XL U8014 ( .A(n23382), .B(n23387), .Y(n22463) );
  NOR2X1 U8015 ( .A(n20512), .B(n20473), .Y(n20520) );
  INVX1 U8016 ( .A(n23227), .Y(n4767) );
  ADDFHX1 U8017 ( .A(n24342), .B(n3069), .CI(n20124), .CO(n20123), .S(n24340)
         );
  NOR2X1 U8018 ( .A(n22378), .B(n23344), .Y(n23337) );
  NOR2X1 U8019 ( .A(n15766), .B(n15765), .Y(n15839) );
  NOR2XL U8020 ( .A(n20568), .B(n20473), .Y(n20465) );
  NOR2XL U8021 ( .A(n9035), .B(n8984), .Y(n8982) );
  NOR2X1 U8022 ( .A(n20508), .B(n20473), .Y(n20395) );
  NOR3X1 U8023 ( .A(n23845), .B(n9035), .C(n8984), .Y(n8991) );
  NAND2X1 U8024 ( .A(n22408), .B(n23237), .Y(n23244) );
  NOR2X1 U8025 ( .A(n22407), .B(n23250), .Y(n23237) );
  NOR2X1 U8026 ( .A(n22377), .B(n22376), .Y(n23322) );
  NAND2X1 U8027 ( .A(n5599), .B(n3515), .Y(n2578) );
  NOR2X1 U8028 ( .A(n22366), .B(n22365), .Y(n23316) );
  NAND2BXL U8029 ( .AN(n20125), .B(n25343), .Y(n25346) );
  NOR2X1 U8030 ( .A(n20447), .B(n20446), .Y(n20476) );
  AOI21X1 U8031 ( .A0(n9028), .A1(n3067), .B0(n9010), .Y(n20477) );
  AOI2BB1X1 U8032 ( .A0N(n22124), .A1N(n22390), .B0(n6188), .Y(n23265) );
  NOR2X1 U8033 ( .A(n22388), .B(n22387), .Y(n23242) );
  OAI21XL U8034 ( .A0(n24868), .A1(n3121), .B0(n23943), .Y(n2580) );
  OR2XL U8035 ( .A(n25269), .B(n25008), .Y(n25009) );
  NOR2X1 U8036 ( .A(n3067), .B(n8953), .Y(n9010) );
  NAND2BXL U8037 ( .AN(n25269), .B(n25268), .Y(n25274) );
  NOR2X1 U8038 ( .A(n22358), .B(n22357), .Y(n23350) );
  NAND2X1 U8039 ( .A(n22271), .B(n22461), .Y(n22199) );
  AOI222XL U8040 ( .A0(n25697), .A1(n20890), .B0(n25743), .B1(y20[31]), .C0(
        n25737), .C1(n25691), .Y(n2391) );
  OR2XL U8041 ( .A(n22385), .B(n3082), .Y(n22346) );
  OAI2BB1XL U8042 ( .A0N(n25728), .A1N(n25727), .B0(n25726), .Y(n25729) );
  XOR2X1 U8043 ( .A(n23412), .B(n22174), .Y(n23411) );
  OR2X1 U8044 ( .A(n20301), .B(n5598), .Y(n5597) );
  NOR2BXL U8045 ( .AN(n22173), .B(n23397), .Y(n22172) );
  OAI21XL U8046 ( .A0(n24843), .A1(n3121), .B0(n23547), .Y(n2582) );
  AOI2BB1X1 U8047 ( .A0N(n22401), .A1N(n22400), .B0(n22399), .Y(n23275) );
  NOR2XL U8048 ( .A(n23393), .B(n22176), .Y(n22174) );
  NAND2BXL U8049 ( .AN(n23546), .B(n4820), .Y(n4819) );
  AND2XL U8050 ( .A(n20725), .B(n20724), .Y(n20720) );
  OAI21XL U8051 ( .A0(n24735), .A1(n3121), .B0(n23938), .Y(n2588) );
  OR2X2 U8052 ( .A(n3031), .B(n9011), .Y(n9007) );
  NOR2X1 U8053 ( .A(n22310), .B(n22309), .Y(n22397) );
  NOR2X1 U8054 ( .A(n22197), .B(n22196), .Y(n22396) );
  INVXL U8055 ( .A(n20095), .Y(n20097) );
  OAI2BB1XL U8056 ( .A0N(n25807), .A1N(n11478), .B0(n5101), .Y(n2604) );
  NAND3BX1 U8057 ( .AN(n3316), .B(n25640), .C(n25639), .Y(n2617) );
  NAND3XL U8058 ( .A(n23564), .B(n23563), .C(n4346), .Y(n2615) );
  OAI21XL U8059 ( .A0(n24582), .A1(n3121), .B0(n23924), .Y(n2602) );
  OR2X2 U8060 ( .A(n3072), .B(n20153), .Y(n20150) );
  NAND2BXL U8061 ( .AN(n23791), .B(n23790), .Y(n5561) );
  OAI21XL U8062 ( .A0(n25594), .A1(n3121), .B0(n23731), .Y(n2610) );
  NAND2BXL U8063 ( .AN(n23936), .B(n23935), .Y(n23937) );
  NAND2X1 U8064 ( .A(n19072), .B(n4345), .Y(n4344) );
  OAI21XL U8065 ( .A0(n4081), .A1(n3121), .B0(n5915), .Y(n2595) );
  INVX4 U8066 ( .A(n20597), .Y(n20576) );
  NOR2BXL U8067 ( .AN(n25644), .B(n4582), .Y(n3316) );
  AND2X1 U8068 ( .A(n23168), .B(n15734), .Y(n23962) );
  NAND2XL U8069 ( .A(n4952), .B(n4970), .Y(n2552) );
  INVXL U8070 ( .A(n23719), .Y(n5356) );
  NAND2BXL U8071 ( .AN(n20774), .B(n4824), .Y(n4823) );
  OAI2BB1XL U8072 ( .A0N(n24319), .A1N(n3065), .B0(n20660), .Y(n2571) );
  OAI21XL U8073 ( .A0(n20691), .A1(n3121), .B0(n5341), .Y(n2534) );
  OAI21X2 U8074 ( .A0(n20790), .A1(n24386), .B0(n5351), .Y(n24319) );
  NAND3X1 U8075 ( .A(n4978), .B(n4975), .C(n4713), .Y(n2543) );
  BUFX3 U8076 ( .A(n24894), .Y(n20182) );
  OAI21XL U8077 ( .A0(n25851), .A1(n4581), .B0(n25130), .Y(n2557) );
  NAND2BXL U8078 ( .AN(n23901), .B(n4846), .Y(n4845) );
  OAI21XL U8079 ( .A0(n3121), .A1(n21029), .B0(n4992), .Y(n2548) );
  NAND2BXL U8080 ( .AN(n23922), .B(n23921), .Y(n23923) );
  NAND2BXL U8081 ( .AN(n20964), .B(n4841), .Y(n4840) );
  NAND2X2 U8082 ( .A(n4348), .B(n4347), .Y(n19072) );
  NAND2BXL U8083 ( .AN(n23473), .B(n23472), .Y(n23474) );
  NAND2BXL U8084 ( .AN(n23507), .B(n23506), .Y(n23508) );
  INVXL U8085 ( .A(n24697), .Y(n24706) );
  NAND3X1 U8086 ( .A(n3460), .B(n3459), .C(n3458), .Y(n2546) );
  AOI21X1 U8087 ( .A0(n4811), .A1(n4579), .B0(n4971), .Y(n4970) );
  NAND2BXL U8088 ( .AN(n11477), .B(n5103), .Y(n5102) );
  NAND2BXL U8089 ( .AN(n23930), .B(n4844), .Y(n4843) );
  AOI21X1 U8090 ( .A0(n20118), .A1(n20117), .B0(n20116), .Y(n20144) );
  NAND2X2 U8091 ( .A(n5010), .B(n5002), .Y(n20712) );
  INVXL U8092 ( .A(n25755), .Y(n25749) );
  INVXL U8093 ( .A(n24888), .Y(n24912) );
  NOR2XL U8094 ( .A(n3973), .B(n24240), .Y(n2282) );
  NAND2BXL U8095 ( .AN(n22188), .B(n22258), .Y(n22260) );
  AOI21XL U8096 ( .A0(n5246), .A1(n25754), .B0(n4255), .Y(n2301) );
  OAI2BB1XL U8097 ( .A0N(n24396), .A1N(n3065), .B0(n24379), .Y(n2526) );
  OAI2BB1XL U8098 ( .A0N(n25199), .A1N(n3065), .B0(n24090), .Y(n2530) );
  OR2X2 U8099 ( .A(n22426), .B(n22193), .Y(n22194) );
  NAND2X1 U8100 ( .A(n4172), .B(n25771), .Y(n25772) );
  OAI2BB1XL U8101 ( .A0N(n25191), .A1N(n3065), .B0(n24339), .Y(n2529) );
  AOI21XL U8102 ( .A0(n25754), .A1(n24696), .B0(n5270), .Y(n2323) );
  NAND2X1 U8103 ( .A(n4893), .B(n25807), .Y(n6109) );
  OR2X2 U8104 ( .A(n25755), .B(n4584), .Y(n4282) );
  AOI22XL U8105 ( .A0(n25195), .A1(n25807), .B0(n2984), .B1(temp1[25]), .Y(
        n24339) );
  AOI22XL U8106 ( .A0(n25204), .A1(n25807), .B0(n2983), .B1(temp1[24]), .Y(
        n24090) );
  AOI22XL U8107 ( .A0(n25166), .A1(n25807), .B0(n2984), .B1(temp1[28]), .Y(
        n24379) );
  INVX1 U8108 ( .A(n3833), .Y(n3832) );
  NAND2X1 U8109 ( .A(n4953), .B(n4954), .Y(n3882) );
  AOI21X1 U8110 ( .A0(n15733), .A1(n15732), .B0(n15731), .Y(n15734) );
  AOI22XL U8111 ( .A0(n25174), .A1(n25807), .B0(n2983), .B1(temp1[27]), .Y(
        n24289) );
  AOI22XL U8112 ( .A0(n25797), .A1(n25807), .B0(n2984), .B1(temp1[30]), .Y(
        n25798) );
  AOI22XL U8113 ( .A0(n25814), .A1(n25807), .B0(n2983), .B1(temp1[23]), .Y(
        n25808) );
  AOI211XL U8114 ( .A0(n25329), .A1(n24220), .B0(n24214), .C0(n24213), .Y(
        n2279) );
  AOI21X4 U8115 ( .A0(n20065), .A1(n20064), .B0(n20063), .Y(n20066) );
  OAI2BB1X2 U8116 ( .A0N(n23883), .A1N(n23626), .B0(n4259), .Y(n5246) );
  NAND2X2 U8117 ( .A(n3463), .B(n3462), .Y(n3461) );
  NOR2X1 U8118 ( .A(n24386), .B(n20781), .Y(n20782) );
  NOR2BX2 U8119 ( .AN(n20065), .B(n20063), .Y(n23200) );
  AOI31X1 U8120 ( .A0(n15726), .A1(n15704), .A2(n15729), .B0(n15703), .Y(
        n24917) );
  INVXL U8121 ( .A(n24847), .Y(n24867) );
  OAI2BB1X2 U8122 ( .A0N(n24127), .A1N(n3353), .B0(n3468), .Y(n5408) );
  INVXL U8123 ( .A(n25197), .Y(n3769) );
  OAI21X1 U8124 ( .A0(n25168), .A1(n4772), .B0(n25167), .Y(n25169) );
  NOR2X1 U8125 ( .A(n24386), .B(n20802), .Y(n20803) );
  NOR2XL U8126 ( .A(n24796), .B(n4586), .Y(n4836) );
  NAND2X2 U8127 ( .A(n3999), .B(n3998), .Y(n4893) );
  AOI22X2 U8128 ( .A0(n4267), .A1(n23747), .B0(n4283), .B1(n3081), .Y(n25755)
         );
  NAND2X1 U8129 ( .A(n3972), .B(n3970), .Y(n25770) );
  NOR2BX2 U8130 ( .AN(n15687), .B(n15685), .Y(n15638) );
  AOI21X4 U8131 ( .A0(n15687), .A1(n15686), .B0(n15685), .Y(n15688) );
  NAND4X1 U8132 ( .A(n8977), .B(n8976), .C(n8973), .D(n8979), .Y(n8934) );
  NAND2X1 U8133 ( .A(n8972), .B(n8968), .Y(n8768) );
  NAND2XL U8134 ( .A(n4852), .B(n4851), .Y(n2308) );
  NAND2X1 U8135 ( .A(n23650), .B(n4267), .Y(n5266) );
  AND2X1 U8136 ( .A(n23114), .B(n23113), .Y(n23225) );
  XOR2X2 U8137 ( .A(n20813), .B(n20812), .Y(n23535) );
  NOR3X1 U8138 ( .A(n15780), .B(n15779), .C(n15778), .Y(n15781) );
  NAND2X1 U8139 ( .A(n3081), .B(n23569), .Y(n4291) );
  NAND2XL U8140 ( .A(n5334), .B(n5337), .Y(n2324) );
  XOR2X2 U8141 ( .A(n5519), .B(n20989), .Y(n23462) );
  NAND2X1 U8142 ( .A(n24200), .B(n20353), .Y(n5334) );
  NAND2X1 U8143 ( .A(n5852), .B(n5851), .Y(mul5_out[16]) );
  AOI22XL U8144 ( .A0(n24237), .A1(n23795), .B0(temp1[18]), .B1(n2983), .Y(
        n23714) );
  INVXL U8145 ( .A(n24350), .Y(n25189) );
  INVXL U8146 ( .A(n20087), .Y(n20089) );
  NAND4X1 U8147 ( .A(n20115), .B(n20114), .C(n20111), .D(n20117), .Y(n20063)
         );
  NOR2X1 U8148 ( .A(n20457), .B(n20458), .Y(n8972) );
  NAND2X2 U8149 ( .A(n4191), .B(n3237), .Y(n3236) );
  OR4X2 U8150 ( .A(n20449), .B(n20450), .C(n20453), .D(n20454), .Y(n8948) );
  NOR2X1 U8151 ( .A(n9030), .B(n20402), .Y(n8977) );
  NAND2X1 U8152 ( .A(n20110), .B(n20106), .Y(n19897) );
  NAND2X1 U8153 ( .A(n11471), .B(n11470), .Y(n20728) );
  NOR2X1 U8154 ( .A(n20542), .B(n20543), .Y(n8973) );
  OAI2BB1X2 U8155 ( .A0N(n3938), .A1N(n4902), .B0(n4063), .Y(n17458) );
  NAND2X1 U8156 ( .A(n11471), .B(n11461), .Y(n20717) );
  INVX1 U8157 ( .A(n9030), .Y(n9031) );
  INVX1 U8158 ( .A(n25834), .Y(n25699) );
  NOR2X1 U8159 ( .A(n20404), .B(n20400), .Y(n8979) );
  XOR2X2 U8160 ( .A(n3666), .B(n2999), .Y(n24192) );
  INVXL U8161 ( .A(n24237), .Y(n4009) );
  NOR3X1 U8162 ( .A(n20435), .B(n20436), .C(n8969), .Y(n8945) );
  NOR2X1 U8163 ( .A(n20561), .B(n20562), .Y(n8976) );
  INVXL U8164 ( .A(n24123), .Y(n4927) );
  NOR2X1 U8165 ( .A(n24938), .B(n24889), .Y(n20114) );
  NAND2BX1 U8166 ( .AN(n6130), .B(n6041), .Y(n24350) );
  XNOR2X1 U8167 ( .A(n8718), .B(n8717), .Y(n20449) );
  CLKINVX4 U8168 ( .A(n25331), .Y(n25329) );
  NOR2X1 U8169 ( .A(n20167), .B(n25343), .Y(n20115) );
  XOR2X2 U8170 ( .A(n4951), .B(n4944), .Y(n24211) );
  XNOR2X1 U8171 ( .A(n8846), .B(n8845), .Y(n20562) );
  XNOR2X1 U8172 ( .A(n8727), .B(n8726), .Y(n20450) );
  XNOR2X1 U8173 ( .A(n8868), .B(n8867), .Y(n20543) );
  NAND4X2 U8174 ( .A(n3235), .B(n3234), .C(n5074), .D(n3233), .Y(n3237) );
  XNOR2X1 U8175 ( .A(n8841), .B(n8840), .Y(n20561) );
  XNOR2X1 U8176 ( .A(n8731), .B(n8730), .Y(n20453) );
  AOI21X1 U8177 ( .A0(n11448), .A1(n11447), .B0(n23673), .Y(n11471) );
  XNOR2X1 U8178 ( .A(n8740), .B(n8739), .Y(n20454) );
  XNOR2X1 U8179 ( .A(n8887), .B(n8886), .Y(n20400) );
  XNOR2X1 U8180 ( .A(n8748), .B(n8747), .Y(n20457) );
  OR4X2 U8181 ( .A(n24798), .B(n24716), .C(n24717), .D(n24680), .Y(n20078) );
  NOR2X1 U8182 ( .A(n20415), .B(n20461), .Y(n8968) );
  NOR3X1 U8183 ( .A(n20195), .B(n20196), .C(n20107), .Y(n20075) );
  XNOR2X1 U8184 ( .A(n8836), .B(n8835), .Y(n20402) );
  OAI21XL U8185 ( .A0(mul5_out[30]), .A1(n3111), .B0(n25787), .Y(n2356) );
  CLKINVX8 U8186 ( .A(n5985), .Y(n3131) );
  NAND4X1 U8187 ( .A(n15730), .B(n15729), .C(n15726), .D(n15732), .Y(n15685)
         );
  NAND2X1 U8188 ( .A(n15725), .B(n15721), .Y(n15517) );
  NAND2X1 U8189 ( .A(n24048), .B(n25789), .Y(n3972) );
  XOR2X1 U8190 ( .A(n19092), .B(n19093), .Y(n23650) );
  NOR2X1 U8191 ( .A(n24849), .B(n24828), .Y(n20111) );
  BUFX8 U8192 ( .A(n3467), .Y(n3353) );
  CLKINVX3 U8193 ( .A(n20707), .Y(n20610) );
  NAND2X1 U8194 ( .A(n8967), .B(n8965), .Y(n8946) );
  NOR2X1 U8195 ( .A(n25344), .B(n24937), .Y(n20117) );
  XOR2X1 U8196 ( .A(n8914), .B(n8913), .Y(n20435) );
  NOR2X1 U8197 ( .A(n24962), .B(n24870), .Y(n15729) );
  NOR2X1 U8198 ( .A(n20439), .B(n20440), .Y(n8967) );
  NOR2X1 U8199 ( .A(n25270), .B(n25007), .Y(n15732) );
  NOR2X1 U8200 ( .A(n24871), .B(n21000), .Y(n15726) );
  OR4X2 U8201 ( .A(n15920), .B(n15923), .C(n15872), .D(n15873), .Y(n15700) );
  NOR3X1 U8202 ( .A(n15819), .B(n15820), .C(n15722), .Y(n15697) );
  NOR2X1 U8203 ( .A(n15860), .B(n15861), .Y(n15725) );
  XOR2X1 U8204 ( .A(n8882), .B(n8850), .Y(n20542) );
  AND2X2 U8205 ( .A(n3667), .B(n3895), .Y(n3666) );
  XOR2X1 U8206 ( .A(n8863), .B(n8757), .Y(n20415) );
  NAND2X1 U8207 ( .A(n23668), .B(n23667), .Y(n25829) );
  NOR2X1 U8208 ( .A(n15782), .B(n25268), .Y(n15730) );
  OAI2BB1X1 U8209 ( .A0N(n25132), .A1N(n23643), .B0(n25109), .Y(mul5_out[29])
         );
  XOR2X1 U8210 ( .A(n4928), .B(n20316), .Y(n24123) );
  AOI21X1 U8211 ( .A0(n22168), .A1(n22167), .B0(n22166), .Y(n22250) );
  XNOR2X1 U8212 ( .A(n19869), .B(n19868), .Y(n24680) );
  XNOR2X1 U8213 ( .A(n19965), .B(n19964), .Y(n25343) );
  XNOR2X1 U8214 ( .A(n20003), .B(n20002), .Y(n25344) );
  XNOR2X1 U8215 ( .A(n19997), .B(n19996), .Y(n24828) );
  XNOR2X1 U8216 ( .A(n19975), .B(n19974), .Y(n24889) );
  NAND2XL U8217 ( .A(n3895), .B(n21035), .Y(n21036) );
  XNOR2X1 U8218 ( .A(n19970), .B(n19969), .Y(n24938) );
  XNOR2X1 U8219 ( .A(n19860), .B(n19859), .Y(n24717) );
  XNOR2X1 U8220 ( .A(n19856), .B(n19855), .Y(n24716) );
  NOR2X1 U8221 ( .A(n20235), .B(n20236), .Y(n20106) );
  XNOR2X1 U8222 ( .A(n20016), .B(n20015), .Y(n24937) );
  XNOR2X1 U8223 ( .A(n19847), .B(n19846), .Y(n24798) );
  XNOR2X1 U8224 ( .A(n15596), .B(n15595), .Y(n24870) );
  NOR2XL U8225 ( .A(n23531), .B(n23533), .Y(n23494) );
  NOR3X1 U8226 ( .A(n22211), .B(n22210), .C(n22209), .Y(n22212) );
  NOR2X1 U8227 ( .A(n15826), .B(n15827), .Y(n15721) );
  NOR2X1 U8228 ( .A(n20443), .B(n9015), .Y(n8965) );
  INVX4 U8229 ( .A(n3261), .Y(n23489) );
  XNOR2X1 U8230 ( .A(n15497), .B(n15496), .Y(n15860) );
  XOR2X1 U8231 ( .A(n19896), .B(n19895), .Y(n20236) );
  XNOR2X1 U8232 ( .A(n15467), .B(n15466), .Y(n15920) );
  NAND2X2 U8233 ( .A(n5174), .B(n4353), .Y(n20947) );
  XNOR2X1 U8234 ( .A(n15476), .B(n15475), .Y(n15923) );
  XNOR2X1 U8235 ( .A(n15502), .B(n15501), .Y(n15861) );
  NAND2X1 U8236 ( .A(n5358), .B(n5357), .Y(n23972) );
  CLKINVX3 U8237 ( .A(n3895), .Y(n5977) );
  INVXL U8238 ( .A(n23573), .Y(n21035) );
  XNOR2X1 U8239 ( .A(n15618), .B(n15617), .Y(n21000) );
  CLKINVX3 U8240 ( .A(n23744), .Y(n3134) );
  OAI2BB1X1 U8241 ( .A0N(n23868), .A1N(n7880), .B0(n7879), .Y(n24447) );
  XNOR2X1 U8242 ( .A(n15624), .B(n15623), .Y(n25270) );
  OAI2BB1X1 U8243 ( .A0N(n23868), .A1N(n23852), .B0(n23851), .Y(n25840) );
  AOI21X4 U8244 ( .A0(n22123), .A1(n22122), .B0(n22121), .Y(n22124) );
  BUFX12 U8245 ( .A(n5335), .Y(n3136) );
  XNOR2X1 U8246 ( .A(n15489), .B(n15488), .Y(n15873) );
  XOR2X1 U8247 ( .A(n17429), .B(n17431), .Y(n17436) );
  XOR2X1 U8248 ( .A(n20011), .B(n19979), .Y(n24849) );
  XNOR2X1 U8249 ( .A(n15579), .B(n15364), .Y(n15782) );
  NOR2XL U8250 ( .A(n5403), .B(n13024), .Y(n5969) );
  NOR2BX2 U8251 ( .AN(n22123), .B(n22121), .Y(n23113) );
  XNOR2X1 U8252 ( .A(n15586), .B(n15585), .Y(n25268) );
  NAND2X1 U8253 ( .A(n20706), .B(n20705), .Y(n20708) );
  INVXL U8254 ( .A(n15872), .Y(n3138) );
  INVXL U8255 ( .A(n20609), .Y(n20706) );
  NAND4X1 U8256 ( .A(n20988), .B(n19074), .C(n4331), .D(n4330), .Y(n10288) );
  OR2XL U8257 ( .A(n15825), .B(n4453), .Y(n15773) );
  XOR2X1 U8258 ( .A(n15632), .B(n15600), .Y(n24871) );
  NAND2X1 U8259 ( .A(n11399), .B(n11470), .Y(n11412) );
  CLKINVX3 U8260 ( .A(n6142), .Y(n5216) );
  AND2X2 U8261 ( .A(n6142), .B(n20636), .Y(n4587) );
  NAND2X1 U8262 ( .A(n3450), .B(n4842), .Y(n24035) );
  NAND3BX2 U8263 ( .AN(n23491), .B(n5317), .C(n5319), .Y(n3261) );
  INVXL U8264 ( .A(n24057), .Y(n4257) );
  XOR2X1 U8265 ( .A(n15613), .B(n15506), .Y(n15826) );
  XOR2X1 U8266 ( .A(n15516), .B(n15515), .Y(n15827) );
  NAND2X2 U8267 ( .A(n20678), .B(n23482), .Y(n4158) );
  NOR2X1 U8268 ( .A(n15835), .B(n15836), .Y(n15718) );
  NAND2BXL U8269 ( .AN(n20269), .B(n4305), .Y(n20609) );
  AND2XL U8270 ( .A(n6198), .B(n23482), .Y(n6199) );
  INVX1 U8271 ( .A(n10226), .Y(n4330) );
  XOR2X2 U8272 ( .A(n5643), .B(n20919), .Y(n20938) );
  XOR2X1 U8273 ( .A(n20352), .B(n20351), .Y(n20943) );
  NAND2BXL U8274 ( .AN(n5569), .B(n23685), .Y(n5571) );
  NAND3X1 U8275 ( .A(n20623), .B(n20286), .C(n11385), .Y(n11399) );
  INVX1 U8276 ( .A(n4306), .Y(n20812) );
  INVXL U8277 ( .A(n23863), .Y(n5568) );
  NAND2XL U8278 ( .A(n5389), .B(n14519), .Y(n14549) );
  NAND4X1 U8279 ( .A(n22165), .B(n22164), .C(n22161), .D(n22167), .Y(n22121)
         );
  XOR2X1 U8280 ( .A(n15647), .B(n15646), .Y(n15825) );
  INVXL U8281 ( .A(n3393), .Y(n17422) );
  CLKINVX3 U8282 ( .A(n3372), .Y(n3374) );
  INVXL U8283 ( .A(n20714), .Y(n20715) );
  XNOR2X1 U8284 ( .A(n8941), .B(n8940), .Y(n9016) );
  INVXL U8285 ( .A(n5389), .Y(n14725) );
  NOR2X1 U8286 ( .A(n5318), .B(n5316), .Y(n23492) );
  NOR2X2 U8287 ( .A(n19048), .B(n4442), .Y(n5228) );
  NAND3X2 U8288 ( .A(n3806), .B(n3627), .C(n5700), .Y(n3373) );
  NAND2X1 U8289 ( .A(n22160), .B(n22156), .Y(n21957) );
  NAND2BXL U8290 ( .AN(n18845), .B(n4198), .Y(n5874) );
  NAND2BX1 U8291 ( .AN(n17457), .B(n17456), .Y(n4043) );
  NOR3X2 U8292 ( .A(n14667), .B(n14666), .C(n14665), .Y(n14671) );
  NOR2X1 U8293 ( .A(n8645), .B(n8924), .Y(n8918) );
  AOI21X2 U8294 ( .A0(n4328), .A1(n10287), .B0(n4326), .Y(n10703) );
  XOR2X1 U8295 ( .A(n17447), .B(n17446), .Y(n20337) );
  XOR2X1 U8296 ( .A(n6045), .B(n20736), .Y(n20935) );
  XOR2X1 U8297 ( .A(n20336), .B(n20335), .Y(n20742) );
  INVXL U8298 ( .A(n6074), .Y(n10709) );
  INVX2 U8299 ( .A(n3911), .Y(n3909) );
  NAND2X2 U8300 ( .A(n3273), .B(n3272), .Y(n20269) );
  OR2XL U8301 ( .A(n23481), .B(n23480), .Y(n6198) );
  INVX1 U8302 ( .A(n4331), .Y(n10713) );
  OR4X2 U8303 ( .A(n22282), .B(n22285), .C(n22286), .D(n22287), .Y(n22136) );
  NOR2X1 U8304 ( .A(n22421), .B(n22252), .Y(n22164) );
  NOR2X1 U8305 ( .A(n22272), .B(n22273), .Y(n22160) );
  INVX1 U8306 ( .A(n15507), .Y(n15680) );
  NAND2X1 U8307 ( .A(n3957), .B(n3357), .Y(n5665) );
  XNOR2X1 U8308 ( .A(n10958), .B(n10957), .Y(n20623) );
  NOR2X1 U8309 ( .A(n22333), .B(n22254), .Y(n22161) );
  XOR2X2 U8310 ( .A(n5588), .B(n20372), .Y(n23807) );
  BUFX2 U8311 ( .A(n20711), .Y(n20713) );
  INVX2 U8312 ( .A(n19074), .Y(n3142) );
  INVX1 U8313 ( .A(n14685), .Y(n20305) );
  AOI21X1 U8314 ( .A0(n15398), .A1(n15667), .B0(n15397), .Y(n15399) );
  NOR2X1 U8315 ( .A(n8774), .B(n8780), .Y(n8784) );
  NOR2X1 U8316 ( .A(n22247), .B(n22244), .Y(n22156) );
  XOR2X2 U8317 ( .A(n5227), .B(n4607), .Y(n20808) );
  XNOR2X1 U8318 ( .A(n22017), .B(n21527), .Y(n22213) );
  NOR2X2 U8319 ( .A(n23651), .B(n20312), .Y(n20670) );
  XNOR2X1 U8320 ( .A(n21916), .B(n21915), .Y(n22285) );
  XNOR2X1 U8321 ( .A(n21942), .B(n21941), .Y(n22273) );
  XNOR2X1 U8322 ( .A(n22024), .B(n22023), .Y(n22258) );
  NOR2X2 U8323 ( .A(n3351), .B(n17359), .Y(n3707) );
  XNOR2X1 U8324 ( .A(n22034), .B(n22033), .Y(n22252) );
  XNOR2X1 U8325 ( .A(n21907), .B(n21906), .Y(n22282) );
  NOR2BX2 U8326 ( .AN(n20371), .B(n4809), .Y(n5588) );
  XNOR2X1 U8327 ( .A(n22029), .B(n22028), .Y(n22421) );
  AND4XL U8328 ( .A(n23541), .B(n20287), .C(n20766), .D(n11384), .Y(n11385) );
  NOR2X1 U8329 ( .A(n5465), .B(n23558), .Y(n5464) );
  XNOR2X1 U8330 ( .A(n21920), .B(n21919), .Y(n22286) );
  NAND3X2 U8331 ( .A(n5409), .B(n2999), .C(n13025), .Y(n3378) );
  OR2XL U8332 ( .A(n23485), .B(n23484), .Y(n6222) );
  AND2X2 U8333 ( .A(n4197), .B(n6032), .Y(n5456) );
  XNOR2X1 U8334 ( .A(n21937), .B(n21936), .Y(n22272) );
  XNOR2X1 U8335 ( .A(n21929), .B(n21928), .Y(n22287) );
  XNOR2X1 U8336 ( .A(n22075), .B(n22074), .Y(n22256) );
  XOR2X1 U8337 ( .A(n22051), .B(n21946), .Y(n22247) );
  NAND2X1 U8338 ( .A(n8851), .B(n8778), .Y(n8780) );
  XNOR2X2 U8339 ( .A(n4329), .B(n10286), .Y(n4328) );
  NAND3X2 U8340 ( .A(n3002), .B(n17470), .C(n3338), .Y(n3351) );
  NAND2X2 U8341 ( .A(n13027), .B(n21043), .Y(n4077) );
  XOR2X1 U8342 ( .A(n22070), .B(n22038), .Y(n22333) );
  NAND4X2 U8343 ( .A(n19044), .B(n5899), .C(n19021), .D(n19020), .Y(n3441) );
  NOR2X2 U8344 ( .A(n5273), .B(n20983), .Y(n4284) );
  INVX1 U8345 ( .A(n15754), .Y(n23956) );
  AOI21X1 U8346 ( .A0(n10971), .A1(n10956), .B0(n10955), .Y(n10961) );
  NOR2XL U8347 ( .A(n20333), .B(n20335), .Y(n17444) );
  CLKINVX3 U8348 ( .A(n20697), .Y(n3445) );
  NOR2X2 U8349 ( .A(n4965), .B(n5410), .Y(n5409) );
  NAND2X2 U8350 ( .A(n2991), .B(n23512), .Y(n4203) );
  NAND3X1 U8351 ( .A(n3596), .B(n5100), .C(n20757), .Y(n20818) );
  INVX1 U8352 ( .A(n13028), .Y(n23572) );
  NOR2X1 U8353 ( .A(n19773), .B(n20053), .Y(n20047) );
  NAND2X1 U8354 ( .A(n3317), .B(n10577), .Y(n10597) );
  NAND2XL U8355 ( .A(n15208), .B(n15649), .Y(n15650) );
  NOR2X2 U8356 ( .A(n4827), .B(n6111), .Y(n6110) );
  INVXL U8357 ( .A(n3956), .Y(n20358) );
  AND2XL U8358 ( .A(n24262), .B(n24261), .Y(n6221) );
  NOR2X1 U8359 ( .A(n8639), .B(n8638), .Y(n8927) );
  AND2X2 U8360 ( .A(n5365), .B(n14544), .Y(n5484) );
  XNOR2X1 U8361 ( .A(n20074), .B(n20073), .Y(n24063) );
  NOR2X1 U8362 ( .A(n8719), .B(n8723), .Y(n8851) );
  NOR2X1 U8363 ( .A(n19903), .B(n19909), .Y(n19913) );
  INVXL U8364 ( .A(n5919), .Y(n5475) );
  NOR2X1 U8365 ( .A(n15523), .B(n15529), .Y(n15533) );
  AOI21X1 U8366 ( .A0(n8819), .A1(n8879), .B0(n8818), .Y(n8869) );
  NAND2X1 U8367 ( .A(n8875), .B(n8819), .Y(n8870) );
  INVX1 U8368 ( .A(n21019), .Y(n21020) );
  NAND2X1 U8369 ( .A(n8741), .B(n8702), .Y(n8774) );
  INVX1 U8370 ( .A(n8523), .Y(n9000) );
  AND2XL U8371 ( .A(n20954), .B(n20953), .Y(n20955) );
  INVX4 U8372 ( .A(n18978), .Y(n3147) );
  AND2XL U8373 ( .A(n20960), .B(n20959), .Y(n20961) );
  AND2XL U8374 ( .A(n15758), .B(n15759), .Y(n15763) );
  NAND3X2 U8375 ( .A(n3956), .B(n20348), .C(n17467), .Y(n3958) );
  AND2X2 U8376 ( .A(n5486), .B(n14536), .Y(n5485) );
  AOI2BB2X2 U8377 ( .B0(n14351), .B1(n4677), .A0N(n14352), .A1N(n4938), .Y(
        n4253) );
  AND2X2 U8378 ( .A(n3326), .B(n10652), .Y(n10654) );
  AND2XL U8379 ( .A(n20146), .B(n20147), .Y(n20151) );
  NAND2X1 U8380 ( .A(n10635), .B(n10638), .Y(n3304) );
  AOI21X1 U8381 ( .A0(n15451), .A1(n15491), .B0(n15450), .Y(n15530) );
  NOR2X1 U8382 ( .A(n8919), .B(n8763), .Y(n8651) );
  NAND2X2 U8383 ( .A(n23458), .B(n23456), .Y(n4404) );
  NOR2BX2 U8384 ( .AN(n12903), .B(n3349), .Y(n3348) );
  NAND2X1 U8385 ( .A(n19980), .B(n19907), .Y(n19909) );
  NOR2BX2 U8386 ( .AN(n12920), .B(n3347), .Y(n3346) );
  NAND2XL U8387 ( .A(n10634), .B(n10588), .Y(n10590) );
  NOR2X1 U8388 ( .A(n8847), .B(n8842), .Y(n8875) );
  NOR2X1 U8389 ( .A(n8856), .B(n8864), .Y(n8778) );
  NAND2X1 U8390 ( .A(n15490), .B(n15451), .Y(n15523) );
  NAND2BX1 U8391 ( .AN(n14352), .B(n3327), .Y(n4939) );
  NOR2X1 U8392 ( .A(n8754), .B(n8749), .Y(n8741) );
  AOI21X1 U8393 ( .A0(n15569), .A1(n15629), .B0(n15568), .Y(n15619) );
  NAND2X1 U8394 ( .A(n15625), .B(n15569), .Y(n15620) );
  BUFX3 U8395 ( .A(n13036), .Y(n4986) );
  OAI21X2 U8396 ( .A0(n3415), .A1(n12869), .B0(n4123), .Y(n4377) );
  NAND2X1 U8397 ( .A(n15601), .B(n15527), .Y(n15529) );
  NOR2X1 U8398 ( .A(n19848), .B(n19852), .Y(n19980) );
  OR2X2 U8399 ( .A(n15369), .B(n15368), .Y(n15261) );
  NOR2X1 U8400 ( .A(n8813), .B(n8812), .Y(n8842) );
  NAND2X1 U8401 ( .A(n8811), .B(n8810), .Y(n8848) );
  NOR2X1 U8402 ( .A(n8706), .B(n8705), .Y(n8723) );
  NOR2X2 U8403 ( .A(n3469), .B(n4647), .Y(n4003) );
  INVX1 U8404 ( .A(n19614), .Y(n20141) );
  NOR2X1 U8405 ( .A(n8715), .B(n8714), .Y(n8856) );
  NAND2X1 U8406 ( .A(n19870), .B(n19831), .Y(n19903) );
  NOR2X1 U8407 ( .A(n8776), .B(n8775), .Y(n8864) );
  NOR2X1 U8408 ( .A(n8696), .B(n8695), .Y(n8749) );
  NOR2X1 U8409 ( .A(n8649), .B(n8648), .Y(n8763) );
  OAI22X1 U8410 ( .A0(n23481), .A1(n14475), .B0(n14474), .B1(n14473), .Y(
        n14662) );
  INVX1 U8411 ( .A(n15274), .Y(n15755) );
  NOR2X1 U8412 ( .A(n15503), .B(n15498), .Y(n15490) );
  OR2XL U8413 ( .A(n23955), .B(n15757), .Y(n15758) );
  NOR2X1 U8414 ( .A(n15669), .B(n15512), .Y(n15398) );
  INVX1 U8415 ( .A(n20739), .Y(n20740) );
  NOR2X1 U8416 ( .A(n15468), .B(n15472), .Y(n15601) );
  NAND3X2 U8417 ( .A(n3525), .B(n3013), .C(n20363), .Y(n3523) );
  NOR2X1 U8418 ( .A(n15606), .B(n15614), .Y(n15527) );
  NOR2X1 U8419 ( .A(n8647), .B(n8646), .Y(n8919) );
  OR2X2 U8420 ( .A(n15376), .B(n15375), .Y(n15208) );
  NOR2X1 U8421 ( .A(n19985), .B(n19993), .Y(n19907) );
  NOR2X1 U8422 ( .A(n8694), .B(n8693), .Y(n8754) );
  NAND2X1 U8423 ( .A(n20004), .B(n19948), .Y(n19999) );
  NOR2X1 U8424 ( .A(n15597), .B(n15592), .Y(n15625) );
  NAND2X1 U8425 ( .A(n4012), .B(n12927), .Y(n4011) );
  NOR2X1 U8426 ( .A(n8811), .B(n8810), .Y(n8847) );
  NOR2X1 U8427 ( .A(n15396), .B(n15395), .Y(n15512) );
  NAND2X2 U8428 ( .A(n20282), .B(n20757), .Y(n3519) );
  NOR2X1 U8429 ( .A(n19844), .B(n19843), .Y(n19985) );
  NAND2X1 U8430 ( .A(n15561), .B(n15560), .Y(n15598) );
  NOR2X1 U8431 ( .A(n19976), .B(n19971), .Y(n20004) );
  NOR2X1 U8432 ( .A(n15561), .B(n15560), .Y(n15597) );
  NOR2X1 U8433 ( .A(n15563), .B(n15562), .Y(n15592) );
  NOR2X1 U8434 ( .A(n19905), .B(n19904), .Y(n19993) );
  NOR2BX2 U8435 ( .AN(n17346), .B(n3793), .Y(n5659) );
  NOR2X1 U8436 ( .A(n8821), .B(n8820), .Y(n8830) );
  NOR2X1 U8437 ( .A(n19775), .B(n19774), .Y(n20048) );
  NOR2X1 U8438 ( .A(n8817), .B(n8816), .Y(n8883) );
  NOR2X1 U8439 ( .A(n15445), .B(n15444), .Y(n15498) );
  NOR2X1 U8440 ( .A(n15525), .B(n15524), .Y(n15614) );
  NOR2X1 U8441 ( .A(n15449), .B(n15448), .Y(n15485) );
  NOR2X1 U8442 ( .A(n19883), .B(n19878), .Y(n19870) );
  NOR2X1 U8443 ( .A(n15443), .B(n15442), .Y(n15503) );
  XNOR2X1 U8444 ( .A(n15348), .B(n15364), .Y(n15757) );
  NOR2X1 U8445 ( .A(n15455), .B(n15454), .Y(n15472) );
  NOR2X1 U8446 ( .A(n15453), .B(n15452), .Y(n15468) );
  NOR2X1 U8447 ( .A(n15571), .B(n15570), .Y(n15580) );
  INVX1 U8448 ( .A(n22185), .Y(n23223) );
  INVX1 U8449 ( .A(n17443), .Y(n20335) );
  INVXL U8450 ( .A(n20365), .Y(n5585) );
  NAND2X1 U8451 ( .A(n7452), .B(n20759), .Y(n3528) );
  NOR2X1 U8452 ( .A(n15394), .B(n15393), .Y(n15669) );
  NAND2X2 U8453 ( .A(n14476), .B(n5150), .Y(n5279) );
  OR2XL U8454 ( .A(n19952), .B(n20145), .Y(n20146) );
  NOR2X1 U8455 ( .A(n15567), .B(n15566), .Y(n15633) );
  INVX1 U8456 ( .A(n14308), .Y(n14352) );
  NOR2BX2 U8457 ( .AN(n10505), .B(n10608), .Y(n4625) );
  NOR2X1 U8458 ( .A(n14351), .B(n4677), .Y(n4263) );
  NOR2X1 U8459 ( .A(n8700), .B(n8699), .Y(n8736) );
  AOI21XL U8460 ( .A0(n10234), .A1(n10233), .B0(n10232), .Y(n10235) );
  INVX1 U8461 ( .A(n20757), .Y(n20815) );
  NAND2X1 U8462 ( .A(n4484), .B(n4482), .Y(n4481) );
  NOR2X1 U8463 ( .A(n14532), .B(n14350), .Y(n14308) );
  NAND2X2 U8464 ( .A(n3604), .B(n5602), .Y(n19060) );
  INVXL U8465 ( .A(n6066), .Y(n14630) );
  NAND3X2 U8466 ( .A(n9762), .B(n3247), .C(n4325), .Y(n3246) );
  NAND2X2 U8467 ( .A(n3247), .B(n4325), .Y(n3244) );
  INVX1 U8468 ( .A(n20363), .Y(n20616) );
  NOR2X1 U8469 ( .A(n19942), .B(n19941), .Y(n19971) );
  NOR2X1 U8470 ( .A(n19940), .B(n19939), .Y(n19976) );
  INVX2 U8471 ( .A(n10182), .Y(n10233) );
  INVXL U8472 ( .A(n17413), .Y(n3850) );
  NOR2X1 U8473 ( .A(n19835), .B(n19834), .Y(n19852) );
  NOR2X1 U8474 ( .A(n19825), .B(n19824), .Y(n19878) );
  NAND3X2 U8475 ( .A(n20816), .B(n20372), .C(n20283), .Y(n3522) );
  NOR2X2 U8476 ( .A(n3242), .B(n3241), .Y(n3240) );
  NAND2X1 U8477 ( .A(n20643), .B(n25241), .Y(n20644) );
  INVX1 U8478 ( .A(n11461), .Y(n11470) );
  AOI2BB1X2 U8479 ( .A0N(n17305), .A1N(n17298), .B0(n4150), .Y(n3960) );
  NOR2X1 U8480 ( .A(n21963), .B(n21969), .Y(n21973) );
  NAND3X2 U8481 ( .A(n4258), .B(n14398), .C(n13982), .Y(n4861) );
  NOR2X1 U8482 ( .A(n19946), .B(n19945), .Y(n20012) );
  AND2X2 U8483 ( .A(n10203), .B(n10202), .Y(n4616) );
  CLKINVX3 U8484 ( .A(n20832), .Y(n3148) );
  AND2XL U8485 ( .A(n11462), .B(n20957), .Y(n11455) );
  INVXL U8486 ( .A(n14483), .Y(n5497) );
  NOR2X1 U8487 ( .A(n19829), .B(n19828), .Y(n19865) );
  XOR2X1 U8488 ( .A(n11398), .B(n11397), .Y(n11461) );
  NOR2X1 U8489 ( .A(n19950), .B(n19949), .Y(n19959) );
  NAND2X1 U8490 ( .A(n15046), .B(n15572), .Y(n15575) );
  OAI2BB1X2 U8491 ( .A0N(n13468), .A1N(n13469), .B0(n5159), .Y(n4258) );
  NAND2X1 U8492 ( .A(n21930), .B(n21891), .Y(n21963) );
  AOI211XL U8493 ( .A0(n9197), .A1(n20790), .B0(n9196), .C0(n20637), .Y(n10666) );
  NAND2X1 U8494 ( .A(n8295), .B(n8822), .Y(n8825) );
  AOI21X1 U8495 ( .A0(n22008), .A1(n22067), .B0(n22007), .Y(n22057) );
  NAND2X1 U8496 ( .A(n22063), .B(n22008), .Y(n22058) );
  NAND2X1 U8497 ( .A(n10646), .B(n10650), .Y(n10653) );
  INVX1 U8498 ( .A(n19076), .Y(n19058) );
  NAND2X1 U8499 ( .A(n8295), .B(n8805), .Y(n8807) );
  NAND2X1 U8500 ( .A(n15046), .B(n15554), .Y(n15556) );
  INVXL U8501 ( .A(n5685), .Y(n5681) );
  INVXL U8502 ( .A(n14636), .Y(n5093) );
  AND2X2 U8503 ( .A(n18915), .B(n18914), .Y(n18916) );
  NAND2X2 U8504 ( .A(n12835), .B(n12780), .Y(n4034) );
  INVX1 U8505 ( .A(n24259), .Y(n3919) );
  NAND2X1 U8506 ( .A(n22039), .B(n21967), .Y(n21969) );
  NAND2X1 U8507 ( .A(n8295), .B(n8800), .Y(n8802) );
  NOR2BX2 U8508 ( .AN(n7427), .B(n3589), .Y(n3588) );
  AOI21X1 U8509 ( .A0(n21891), .A1(n21931), .B0(n21890), .Y(n21970) );
  NOR2X1 U8510 ( .A(n10056), .B(n10055), .Y(n3248) );
  NAND2BXL U8511 ( .AN(n17371), .B(n17390), .Y(n5685) );
  NOR2X2 U8512 ( .A(n4324), .B(n5138), .Y(n3243) );
  ADDFHX2 U8513 ( .A(n10116), .B(n10114), .CI(n10115), .CO(n10117), .S(n10058)
         );
  NAND3BX1 U8514 ( .AN(n7434), .B(n4545), .C(n4544), .Y(n4543) );
  NOR2X1 U8515 ( .A(n10585), .B(n10591), .Y(n10646) );
  XOR2X2 U8516 ( .A(n7017), .B(n7016), .Y(n5602) );
  NAND2X2 U8517 ( .A(n14556), .B(n14570), .Y(n14521) );
  NOR2X1 U8518 ( .A(n22106), .B(n21952), .Y(n21836) );
  AOI21X2 U8519 ( .A0(n10050), .A1(n3256), .B0(n10049), .Y(n3255) );
  INVXL U8520 ( .A(n14551), .Y(n14569) );
  NOR2X2 U8521 ( .A(n14312), .B(n14311), .Y(n14573) );
  NOR2X1 U8522 ( .A(n21908), .B(n21912), .Y(n22039) );
  NOR2X1 U8523 ( .A(n22044), .B(n22052), .Y(n21967) );
  NAND2X2 U8524 ( .A(n13983), .B(n13984), .Y(n14636) );
  NAND2X2 U8525 ( .A(n5367), .B(n12419), .Y(n3714) );
  NAND2X2 U8526 ( .A(n13993), .B(n13992), .Y(n14625) );
  NOR2X1 U8527 ( .A(n21943), .B(n21938), .Y(n21930) );
  NOR2X2 U8528 ( .A(n17225), .B(n3366), .Y(n3365) );
  NOR2X1 U8529 ( .A(n22035), .B(n22030), .Y(n22063) );
  NAND2X2 U8530 ( .A(n3254), .B(n3250), .Y(n3249) );
  NAND2X2 U8531 ( .A(n10131), .B(n10130), .Y(n10220) );
  NAND2X1 U8532 ( .A(n3087), .B(n8437), .Y(n8511) );
  NOR2X1 U8533 ( .A(n21883), .B(n21882), .Y(n21943) );
  NOR2X4 U8534 ( .A(n8614), .B(n8610), .Y(n8295) );
  NAND2BX1 U8535 ( .AN(n20637), .B(n20636), .Y(n20638) );
  NAND2X2 U8536 ( .A(n3089), .B(n3088), .Y(n14570) );
  AND2X2 U8537 ( .A(n12888), .B(n12887), .Y(n12889) );
  AND2X2 U8538 ( .A(n12883), .B(n12931), .Y(n12932) );
  NAND2X1 U8539 ( .A(n12899), .B(n12898), .Y(n12900) );
  NAND2X2 U8540 ( .A(n3680), .B(n17206), .Y(n3364) );
  NOR2X1 U8541 ( .A(n15262), .B(n3090), .Y(n15554) );
  AND2X2 U8542 ( .A(n10285), .B(n10284), .Y(n10286) );
  NOR2BX2 U8543 ( .AN(n9833), .B(n9832), .Y(n3254) );
  NOR2X1 U8544 ( .A(n22010), .B(n22009), .Y(n22018) );
  ADDFHX2 U8545 ( .A(n13823), .B(n13822), .CI(n13821), .CO(n13985), .S(n13984)
         );
  AND2X2 U8546 ( .A(n12876), .B(n12875), .Y(n12877) );
  ADDFHX2 U8547 ( .A(n14039), .B(n14038), .CI(n14037), .CO(n14312), .S(n14309)
         );
  NOR2X1 U8548 ( .A(n21889), .B(n21888), .Y(n21925) );
  NAND2X2 U8549 ( .A(n17124), .B(n17312), .Y(n4103) );
  AND2X2 U8550 ( .A(n18911), .B(n18909), .Y(n18908) );
  NOR2X1 U8551 ( .A(n21895), .B(n21894), .Y(n21912) );
  NOR2X1 U8552 ( .A(n22006), .B(n22005), .Y(n22071) );
  INVXL U8553 ( .A(n10206), .Y(n4352) );
  NOR2X1 U8554 ( .A(n21965), .B(n21964), .Y(n22052) );
  NOR2X1 U8555 ( .A(n21834), .B(n21833), .Y(n21952) );
  NAND2X1 U8556 ( .A(n19424), .B(n19951), .Y(n19954) );
  OAI2BB1X2 U8557 ( .A0N(n10040), .A1N(n10041), .B0(n3251), .Y(n3250) );
  ADDFHX2 U8558 ( .A(n9689), .B(n9688), .CI(n9687), .CO(n10057), .S(n10056) );
  NAND2X1 U8559 ( .A(n19424), .B(n19934), .Y(n19936) );
  NOR2X1 U8560 ( .A(n23659), .B(n9187), .Y(n9197) );
  NOR2X1 U8561 ( .A(n22000), .B(n21999), .Y(n22035) );
  INVXL U8562 ( .A(n10574), .Y(n10578) );
  NOR2X1 U8563 ( .A(n22002), .B(n22001), .Y(n22030) );
  ADDFHX2 U8564 ( .A(n9488), .B(n9487), .CI(n9486), .CO(n10136), .S(n10134) );
  NAND2X1 U8565 ( .A(n12983), .B(n12982), .Y(n4624) );
  NOR2X1 U8566 ( .A(n21832), .B(n21831), .Y(n22106) );
  INVX1 U8567 ( .A(n3328), .Y(n17335) );
  OAI21X2 U8568 ( .A0(n3474), .A1(n3473), .B0(n3471), .Y(n12425) );
  ADDFHX2 U8569 ( .A(n9409), .B(n9408), .CI(n9407), .CO(n9371), .S(n9410) );
  OAI2BB1X2 U8570 ( .A0N(n17367), .A1N(n17362), .B0(n17366), .Y(n4107) );
  INVXL U8571 ( .A(n17242), .Y(n17238) );
  AOI21X1 U8572 ( .A0(n12989), .A1(n12988), .B0(n12987), .Y(n12990) );
  XOR2X1 U8573 ( .A(n9763), .B(n3279), .Y(n10054) );
  NOR2X1 U8574 ( .A(n10521), .B(n10556), .Y(n10574) );
  ADDFHX2 U8575 ( .A(n14010), .B(n14009), .CI(n14008), .CO(n14038), .S(n14002)
         );
  INVX1 U8576 ( .A(n19000), .Y(n19001) );
  CLKINVX2 U8577 ( .A(n14315), .Y(n4271) );
  NAND2X2 U8578 ( .A(n3361), .B(n5338), .Y(n3360) );
  XNOR2X1 U8579 ( .A(n20640), .B(n20639), .Y(n20637) );
  INVX1 U8580 ( .A(n3252), .Y(n3251) );
  NAND2X2 U8581 ( .A(n14535), .B(n14337), .Y(n14503) );
  AOI21XL U8582 ( .A0(n17417), .A1(n17416), .B0(n17415), .Y(n17418) );
  OAI21XL U8583 ( .A0(n21854), .A1(n22013), .B0(n22012), .Y(n22023) );
  NOR2X1 U8584 ( .A(n19600), .B(n19807), .Y(n19934) );
  NAND2X1 U8585 ( .A(n17247), .B(n17246), .Y(n17248) );
  NAND2X1 U8586 ( .A(n13826), .B(n13825), .Y(n6046) );
  ADDFHX2 U8587 ( .A(n9418), .B(n9417), .CI(n9416), .CO(n9411), .S(n10060) );
  NAND2X1 U8588 ( .A(n18325), .B(n17985), .Y(n18328) );
  INVX1 U8589 ( .A(n14399), .Y(n3152) );
  ADDFHX2 U8590 ( .A(n13946), .B(n13944), .CI(n13945), .CO(n13999), .S(n13997)
         );
  INVX1 U8591 ( .A(n15278), .Y(n15040) );
  ADDFHX2 U8592 ( .A(n14163), .B(n14162), .CI(n14161), .CO(n14313), .S(n14311)
         );
  ADDFHX2 U8593 ( .A(n9560), .B(n9559), .CI(n9558), .CO(n10143), .S(n10141) );
  ADDFHX2 U8594 ( .A(n9557), .B(n9556), .CI(n9555), .CO(n10140), .S(n10138) );
  INVXL U8595 ( .A(n5176), .Y(n5179) );
  NAND2X1 U8596 ( .A(n7022), .B(n7021), .Y(n7023) );
  NOR2X1 U8597 ( .A(n19688), .B(n19807), .Y(n19951) );
  NAND2X1 U8598 ( .A(n3253), .B(n10037), .Y(n3252) );
  OR2XL U8599 ( .A(n21575), .B(n21787), .Y(n21577) );
  AOI21X1 U8600 ( .A0(n18325), .A1(n18324), .B0(n18323), .Y(n18326) );
  NAND2X1 U8601 ( .A(n18836), .B(n18835), .Y(n18837) );
  NAND2X2 U8602 ( .A(n12779), .B(n12611), .Y(n4056) );
  NAND2X1 U8603 ( .A(n12767), .B(n12768), .Y(n12979) );
  NAND2X1 U8604 ( .A(n12912), .B(n3844), .Y(n12913) );
  AND2X2 U8605 ( .A(n12611), .B(n12856), .Y(n12857) );
  NAND2X1 U8606 ( .A(n5528), .B(n5527), .Y(n10320) );
  NAND2X1 U8607 ( .A(n12984), .B(n12988), .Y(n12991) );
  NAND2X1 U8608 ( .A(n17360), .B(n17367), .Y(n17144) );
  NAND2X1 U8609 ( .A(n12911), .B(n12910), .Y(n4590) );
  INVX1 U8610 ( .A(n12879), .Y(n12880) );
  NOR2X1 U8611 ( .A(n8606), .B(n8372), .Y(n8437) );
  INVXL U8612 ( .A(n10428), .Y(n6164) );
  INVX1 U8613 ( .A(n17312), .Y(n17324) );
  AND2X2 U8614 ( .A(n17297), .B(n17295), .Y(n17228) );
  NOR2X1 U8615 ( .A(n14657), .B(n14656), .Y(n14660) );
  NOR2XL U8616 ( .A(n10551), .B(n10644), .Y(n5257) );
  NOR2X1 U8617 ( .A(n15031), .B(n15030), .Y(n15329) );
  NAND2XL U8618 ( .A(n10043), .B(n10042), .Y(n10045) );
  NAND2X2 U8619 ( .A(n4910), .B(n5961), .Y(n12863) );
  XNOR2X1 U8620 ( .A(n8278), .B(n8277), .Y(n8284) );
  INVXL U8621 ( .A(n10044), .Y(n5178) );
  NAND2X1 U8622 ( .A(n17301), .B(n17300), .Y(n17302) );
  INVXL U8623 ( .A(n6043), .Y(n6042) );
  XNOR2X1 U8624 ( .A(n15039), .B(n6195), .Y(n15278) );
  OAI2BB1XL U8625 ( .A0N(n14111), .A1N(n14110), .B0(n14109), .Y(n14138) );
  ADDFHX2 U8626 ( .A(n14114), .B(n14112), .CI(n14113), .CO(n14137), .S(n14177)
         );
  AOI21X2 U8627 ( .A0(n18694), .A1(n18928), .B0(n18693), .Y(n18984) );
  NAND2X2 U8628 ( .A(n16845), .B(n16844), .Y(n17261) );
  ADDFHX2 U8629 ( .A(n13952), .B(n13951), .CI(n13950), .CO(n14003), .S(n13945)
         );
  ADDFHX2 U8630 ( .A(n9349), .B(n9348), .CI(n9347), .CO(n9487), .S(n9369) );
  NAND2XL U8631 ( .A(n6160), .B(n6159), .Y(n6158) );
  ADDFHX2 U8632 ( .A(n13805), .B(n13804), .CI(n13803), .CO(n13754), .S(n13823)
         );
  NOR2X1 U8633 ( .A(n3035), .B(n19502), .Y(n19714) );
  OAI21X1 U8634 ( .A0(n9692), .A1(n9691), .B0(n9690), .Y(n6068) );
  NOR2XL U8635 ( .A(n13340), .B(n13341), .Y(n4477) );
  ADDFHX2 U8636 ( .A(n13750), .B(n13749), .CI(n13748), .CO(n13756), .S(n13813)
         );
  NAND2X1 U8637 ( .A(n21506), .B(n21994), .Y(n21996) );
  NAND2X1 U8638 ( .A(n14646), .B(n14651), .Y(n14346) );
  NAND2X1 U8639 ( .A(n25241), .B(n25240), .Y(n20646) );
  ADDFHX2 U8640 ( .A(n13589), .B(n13588), .CI(n13587), .CO(n13595), .S(n13593)
         );
  INVX4 U8641 ( .A(n8668), .Y(n3160) );
  XNOR2X2 U8642 ( .A(n13806), .B(n5327), .Y(n13815) );
  NOR2X1 U8643 ( .A(n10482), .B(n10481), .Y(n10521) );
  ADDFHX2 U8644 ( .A(n10101), .B(n10100), .CI(n10099), .CO(n10121), .S(n10120)
         );
  NOR2X1 U8645 ( .A(n10564), .B(n10563), .Y(n10591) );
  NOR2X1 U8646 ( .A(n10560), .B(n10559), .Y(n10582) );
  ADDFHX2 U8647 ( .A(n9352), .B(n9351), .CI(n9350), .CO(n9485), .S(n9348) );
  XOR3X2 U8648 ( .A(n10438), .B(n10439), .C(n10437), .Y(n10429) );
  AOI21X2 U8649 ( .A0(n3514), .A1(n5551), .B0(n5549), .Y(n3513) );
  XNOR2X1 U8650 ( .A(n15029), .B(n15028), .Y(n15030) );
  NAND2X1 U8651 ( .A(n17370), .B(n17139), .Y(n17387) );
  NAND2X2 U8652 ( .A(n5057), .B(n5686), .Y(n17339) );
  OAI21X2 U8653 ( .A0(n3902), .A1(n3898), .B0(n3896), .Y(n11787) );
  NOR2X1 U8654 ( .A(n14506), .B(n14514), .Y(n14646) );
  AOI2BB2X1 U8655 ( .B0(n24027), .B1(n24028), .A0N(n24028), .A1N(n24027), .Y(
        n24025) );
  XNOR2X1 U8656 ( .A(n8286), .B(n8282), .Y(n8283) );
  ADDFHX2 U8657 ( .A(n14169), .B(n14168), .CI(n14167), .CO(n14176), .S(n14174)
         );
  INVX1 U8658 ( .A(n8528), .Y(n8289) );
  AND2X2 U8659 ( .A(n18322), .B(n18321), .Y(n18323) );
  ADDFHX2 U8660 ( .A(n10147), .B(n10146), .CI(n10145), .CO(n10176), .S(n10142)
         );
  INVXL U8661 ( .A(n12844), .Y(n3988) );
  NAND2XL U8662 ( .A(n13198), .B(n13191), .Y(n13200) );
  INVX1 U8663 ( .A(n10038), .Y(n3238) );
  INVXL U8664 ( .A(n12421), .Y(n3712) );
  ADDFHX2 U8665 ( .A(n13524), .B(n13523), .CI(n13522), .CO(n13588), .S(n13547)
         );
  OAI2BB1X2 U8666 ( .A0N(n16805), .A1N(n16804), .B0(n3681), .Y(n16782) );
  OR2X2 U8667 ( .A(n4237), .B(n12384), .Y(n4236) );
  ADDFHX1 U8668 ( .A(n14181), .B(n14180), .CI(n14179), .CO(n14324), .S(n14319)
         );
  NAND2X1 U8669 ( .A(n3615), .B(n3614), .Y(n16777) );
  XNOR2X2 U8670 ( .A(n12687), .B(n6114), .Y(n4073) );
  INVXL U8671 ( .A(n12905), .Y(n4949) );
  XOR2X2 U8672 ( .A(n8294), .B(n8293), .Y(n8610) );
  AOI21XL U8673 ( .A0(n24349), .A1(n4698), .B0(n6133), .Y(n6043) );
  NOR2X1 U8674 ( .A(n10670), .B(n10669), .Y(n25241) );
  XNOR2X1 U8675 ( .A(n15021), .B(n15020), .Y(n15031) );
  INVX1 U8676 ( .A(n17237), .Y(n3161) );
  NOR2X1 U8677 ( .A(n3092), .B(n8553), .Y(n8372) );
  OAI21X2 U8678 ( .A0(n4026), .A1(n4025), .B0(n4024), .Y(n11862) );
  ADDFHX2 U8679 ( .A(n13457), .B(n13456), .CI(n13455), .CO(n13464), .S(n13462)
         );
  INVXL U8680 ( .A(n17646), .Y(n6160) );
  XOR3X2 U8681 ( .A(n17647), .B(n17646), .C(n17645), .Y(n18406) );
  NOR2X1 U8682 ( .A(n19414), .B(n19413), .Y(n19654) );
  XOR2XL U8683 ( .A(n25776), .B(n25775), .Y(n25777) );
  ADDFHX2 U8684 ( .A(n13940), .B(n13939), .CI(n13938), .CO(n13944), .S(n13941)
         );
  ADDFHX2 U8685 ( .A(n12088), .B(n12087), .CI(n12086), .CO(n12427), .S(n12426)
         );
  AND2X2 U8686 ( .A(n18320), .B(n18319), .Y(n18324) );
  NAND2BXL U8687 ( .AN(n17133), .B(n5082), .Y(n5081) );
  AND2X2 U8688 ( .A(n18859), .B(n18858), .Y(n18860) );
  INVXL U8689 ( .A(n13310), .Y(n4262) );
  INVXL U8690 ( .A(n13309), .Y(n4261) );
  ADDFHX1 U8691 ( .A(n9720), .B(n9719), .CI(n9718), .CO(n9716), .S(n9767) );
  NAND2X1 U8692 ( .A(n7814), .B(n7818), .Y(n7821) );
  INVXL U8693 ( .A(n21787), .Y(n21805) );
  XOR2X1 U8694 ( .A(n4018), .B(n12214), .Y(n12416) );
  NAND2X1 U8695 ( .A(n8292), .B(n8291), .Y(n8293) );
  ADDFHX2 U8696 ( .A(n13338), .B(n13337), .CI(n13336), .CO(n13347), .S(n13343)
         );
  ADDFHX2 U8697 ( .A(n13307), .B(n13306), .CI(n13305), .CO(n13342), .S(n13341)
         );
  AND2X2 U8698 ( .A(n18854), .B(n18855), .Y(n18856) );
  ADDFHX2 U8699 ( .A(n9271), .B(n9270), .CI(n9269), .CO(n9349), .S(n9329) );
  NOR2X1 U8700 ( .A(n19006), .B(n19015), .Y(n18992) );
  XOR3X2 U8701 ( .A(n11825), .B(n11824), .C(n11823), .Y(n11864) );
  XNOR2X1 U8702 ( .A(n8288), .B(n6178), .Y(n8528) );
  ADDFHX2 U8703 ( .A(n13419), .B(n13418), .CI(n13417), .CO(n13459), .S(n13348)
         );
  NAND2X1 U8704 ( .A(n18847), .B(n18855), .Y(n18926) );
  AND2X2 U8705 ( .A(n7440), .B(n7439), .Y(n7441) );
  INVX1 U8706 ( .A(n8272), .Y(n8252) );
  INVX1 U8707 ( .A(n18321), .Y(n5506) );
  NOR2X1 U8708 ( .A(n14341), .B(n14340), .Y(n14514) );
  AND2XL U8709 ( .A(n13195), .B(n13194), .Y(n13196) );
  ADDFHX2 U8710 ( .A(n9336), .B(n9335), .CI(n9334), .CO(n9454), .S(n9367) );
  XOR3X2 U8711 ( .A(n12481), .B(n12480), .C(n3908), .Y(n12482) );
  INVX1 U8712 ( .A(n10720), .Y(n10725) );
  INVX4 U8713 ( .A(n19796), .Y(n3165) );
  ADDFHX2 U8714 ( .A(n18358), .B(n18357), .CI(n18356), .CO(n18398), .S(n18397)
         );
  NAND2X1 U8715 ( .A(n16803), .B(n3682), .Y(n3681) );
  XOR2X2 U8716 ( .A(n5664), .B(n17026), .Y(n17106) );
  XNOR2X1 U8717 ( .A(n19408), .B(n19407), .Y(n19414) );
  NAND2XL U8718 ( .A(n14020), .B(n6098), .Y(n6097) );
  OR2X2 U8719 ( .A(n14332), .B(n14331), .Y(n14272) );
  ADDFHX1 U8720 ( .A(n14144), .B(n14143), .CI(n14142), .CO(n14180), .S(n14136)
         );
  NAND2X1 U8721 ( .A(n24049), .B(n24050), .Y(n4500) );
  OR2X2 U8722 ( .A(n12406), .B(n12405), .Y(n4234) );
  ADDFHX2 U8723 ( .A(n17016), .B(n17014), .CI(n17015), .CO(n17107), .S(n16864)
         );
  XOR3X2 U8724 ( .A(n4146), .B(n13979), .C(n13978), .Y(n13948) );
  ADDFHX2 U8725 ( .A(n10378), .B(n10377), .CI(n10376), .CO(n10393), .S(n10425)
         );
  ADDFHX2 U8726 ( .A(n14172), .B(n14171), .CI(n14170), .CO(n14173), .S(n14162)
         );
  ADDFHX2 U8727 ( .A(n13922), .B(n13921), .CI(n13920), .CO(n13951), .S(n13939)
         );
  ADDFHX2 U8728 ( .A(n18334), .B(n18333), .CI(n18332), .CO(n18401), .S(n18399)
         );
  NAND2XL U8729 ( .A(n9830), .B(n9831), .Y(n5743) );
  NAND2XL U8730 ( .A(n10066), .B(n10067), .Y(n4564) );
  OR2X2 U8731 ( .A(n14330), .B(n14329), .Y(n14495) );
  NOR2X1 U8732 ( .A(n7487), .B(n7490), .Y(n7779) );
  XNOR3X2 U8733 ( .A(n12217), .B(n12216), .C(n4004), .Y(n12411) );
  NAND2X1 U8734 ( .A(n7770), .B(n7769), .Y(n4680) );
  INVX1 U8735 ( .A(n19619), .Y(n19418) );
  XNOR2X1 U8736 ( .A(n19406), .B(n19412), .Y(n19413) );
  XNOR2X1 U8737 ( .A(n3997), .B(n12385), .Y(n12406) );
  INVXL U8738 ( .A(n16077), .Y(n6118) );
  NAND2X1 U8739 ( .A(n7668), .B(n7786), .Y(n7670) );
  ADDFHX2 U8740 ( .A(n18388), .B(n18387), .CI(n18386), .CO(n18396), .S(n18395)
         );
  NAND2XL U8741 ( .A(n4355), .B(n4354), .Y(n10420) );
  AND2X2 U8742 ( .A(n23644), .B(n23645), .Y(n5738) );
  OAI2BB1X1 U8743 ( .A0N(n3386), .A1N(n12133), .B0(n3384), .Y(n12111) );
  ADDFHX2 U8744 ( .A(n13765), .B(n13764), .CI(n13763), .CO(n13832), .S(n13761)
         );
  OAI21XL U8745 ( .A0(n4961), .A1(n5792), .B0(n5791), .Y(n12408) );
  OAI21X2 U8746 ( .A0(n5000), .A1(n4999), .B0(n4998), .Y(n12673) );
  ADDFHX2 U8747 ( .A(n18379), .B(n18378), .CI(n18377), .CO(n18390), .S(n18383)
         );
  NAND2BXL U8748 ( .AN(n14021), .B(n6100), .Y(n6098) );
  NAND2BXL U8749 ( .AN(n9519), .B(n5171), .Y(n5170) );
  NOR2X1 U8750 ( .A(n10721), .B(n10722), .Y(n10720) );
  ADDFHX2 U8751 ( .A(n13835), .B(n13834), .CI(n13833), .CO(n13885), .S(n13831)
         );
  ADDFHX2 U8752 ( .A(n13925), .B(n13924), .CI(n13923), .CO(n13949), .S(n13920)
         );
  INVXL U8753 ( .A(n21768), .Y(n21571) );
  AND2X2 U8754 ( .A(n17352), .B(n17351), .Y(n4630) );
  INVXL U8755 ( .A(n4019), .Y(n4017) );
  INVX1 U8756 ( .A(n24046), .Y(n5934) );
  INVXL U8757 ( .A(n20650), .Y(n6032) );
  INVXL U8758 ( .A(n17027), .Y(n5662) );
  NAND2X1 U8759 ( .A(n15043), .B(n15042), .Y(n15044) );
  ADDFHX2 U8760 ( .A(n16452), .B(n16451), .CI(n16450), .CO(n16780), .S(n16779)
         );
  ADDFHX2 U8761 ( .A(n13713), .B(n13712), .CI(n13711), .CO(n13762), .S(n13755)
         );
  INVX1 U8762 ( .A(n12722), .Y(n12977) );
  NAND2BXL U8763 ( .AN(n9825), .B(n5284), .Y(n5283) );
  NAND2BXL U8764 ( .AN(n13501), .B(n4496), .Y(n4495) );
  NOR2XL U8765 ( .A(n12976), .B(n12736), .Y(n5992) );
  AND2X2 U8766 ( .A(n12843), .B(n12842), .Y(n12844) );
  INVX1 U8767 ( .A(n12848), .Y(n12840) );
  AND2X2 U8768 ( .A(n4634), .B(n17358), .Y(n4683) );
  NAND2BXL U8769 ( .AN(n9650), .B(n5196), .Y(n5195) );
  ADDFHX2 U8770 ( .A(n16841), .B(n16840), .CI(n16839), .CO(n16842), .S(n16781)
         );
  NOR2XL U8771 ( .A(n15791), .B(n15790), .Y(n23960) );
  XNOR2X2 U8772 ( .A(n4032), .B(n12678), .Y(n12685) );
  NAND2X1 U8773 ( .A(n9142), .B(n10681), .Y(n9139) );
  OAI2BB1XL U8774 ( .A0N(n9422), .A1N(n5532), .B0(n5531), .Y(n9393) );
  INVXL U8775 ( .A(n5766), .Y(n4557) );
  CLKINVX3 U8776 ( .A(n15128), .Y(n3167) );
  OAI2BB1X1 U8777 ( .A0N(n3267), .A1N(n9376), .B0(n3265), .Y(n9315) );
  NAND2XL U8778 ( .A(n13662), .B(n13661), .Y(n13663) );
  NOR2X2 U8779 ( .A(n18416), .B(n18417), .Y(n18881) );
  AND2X2 U8780 ( .A(n7873), .B(n7872), .Y(n4689) );
  ADDFHX2 U8781 ( .A(n9311), .B(n9310), .CI(n9309), .CO(n9330), .S(n9408) );
  ADDFHX2 U8782 ( .A(n11964), .B(n11963), .CI(n11962), .CO(n12509), .S(n12507)
         );
  XOR2X1 U8783 ( .A(n12215), .B(n4019), .Y(n4018) );
  ADDFHX1 U8784 ( .A(n10070), .B(n10069), .CI(n10068), .CO(n10067), .S(n10098)
         );
  ADDFHX2 U8785 ( .A(n11872), .B(n11871), .CI(n11870), .CO(n11903), .S(n11899)
         );
  XOR2X1 U8786 ( .A(n5261), .B(n13440), .Y(n13437) );
  NAND2X1 U8787 ( .A(n15785), .B(n23966), .Y(n15792) );
  ADDFHX2 U8788 ( .A(n16455), .B(n16454), .CI(n16453), .CO(n16778), .S(n16776)
         );
  AOI21X1 U8789 ( .A0(n15016), .A1(n15015), .B0(n15014), .Y(n15045) );
  XOR3X2 U8790 ( .A(n12432), .B(n12431), .C(n12430), .Y(n12487) );
  INVXL U8791 ( .A(n12386), .Y(n5792) );
  NAND2XL U8792 ( .A(n6052), .B(n23174), .Y(n6051) );
  INVXL U8793 ( .A(n9789), .Y(n5766) );
  NAND2XL U8794 ( .A(n9650), .B(n9649), .Y(n5194) );
  NAND2BXL U8795 ( .AN(n9246), .B(n4309), .Y(n4308) );
  AND2X1 U8796 ( .A(n17393), .B(n17392), .Y(n4692) );
  NAND2XL U8797 ( .A(n9519), .B(n9520), .Y(n5169) );
  NAND2XL U8798 ( .A(n9824), .B(n9825), .Y(n5282) );
  OR2X2 U8799 ( .A(n24431), .B(n15027), .Y(n15026) );
  INVX1 U8800 ( .A(n19401), .Y(n19382) );
  XOR2X1 U8801 ( .A(n9245), .B(n4310), .Y(n9255) );
  ADDFHX2 U8802 ( .A(n18373), .B(n18372), .CI(n18371), .CO(n18357), .S(n18386)
         );
  OAI2BB1XL U8803 ( .A0N(n5242), .A1N(n9247), .B0(n5241), .Y(n9257) );
  INVXL U8804 ( .A(n9520), .Y(n5171) );
  INVXL U8805 ( .A(n17028), .Y(n5663) );
  XOR2X1 U8806 ( .A(n12476), .B(n5775), .Y(n3742) );
  XNOR2X1 U8807 ( .A(n19417), .B(n6200), .Y(n19619) );
  NOR2X1 U8808 ( .A(n9145), .B(n10677), .Y(n9142) );
  INVXL U8809 ( .A(n17351), .Y(n5082) );
  INVXL U8810 ( .A(n5215), .Y(n5214) );
  ADDFHX2 U8811 ( .A(n16823), .B(n16822), .CI(n16821), .CO(n16807), .S(n16824)
         );
  NAND2BX1 U8812 ( .AN(n23634), .B(n23633), .Y(n23635) );
  ADDFHX2 U8813 ( .A(n4748), .B(n9237), .CI(n9236), .CO(n9270), .S(n9310) );
  NOR2X1 U8814 ( .A(n7305), .B(n7304), .Y(n7487) );
  NOR2X1 U8815 ( .A(n7876), .B(n7875), .Y(n10722) );
  ADDFHX2 U8816 ( .A(n10092), .B(n10091), .CI(n10090), .CO(n10085), .S(n10109)
         );
  NOR2X1 U8817 ( .A(n18703), .B(n18942), .Y(n18979) );
  NOR2X1 U8818 ( .A(n16765), .B(n16764), .Y(n16766) );
  INVXL U8819 ( .A(n14021), .Y(n6099) );
  ADDFHX2 U8820 ( .A(n13386), .B(n13385), .CI(n13384), .CO(n13439), .S(n13412)
         );
  ADDFHX2 U8821 ( .A(n13301), .B(n13300), .CI(n13299), .CO(n13306), .S(n13308)
         );
  ADDFHX2 U8822 ( .A(n9429), .B(n9428), .CI(n9427), .CO(n9413), .S(n10066) );
  NAND4X1 U8823 ( .A(n14961), .B(n14960), .C(n14959), .D(n14958), .Y(n14962)
         );
  NOR3X1 U8824 ( .A(n23634), .B(n17265), .C(n17202), .Y(n17394) );
  XOR2X1 U8825 ( .A(n13442), .B(n13441), .Y(n5261) );
  ADDFHX2 U8826 ( .A(n17812), .B(n17810), .CI(n17811), .CO(n18417), .S(n18415)
         );
  NOR2X1 U8827 ( .A(n20374), .B(n8275), .Y(n8279) );
  NAND2BX2 U8828 ( .AN(n6729), .B(n3572), .Y(n6417) );
  XNOR2X1 U8829 ( .A(n14083), .B(n4278), .Y(n4277) );
  NAND2X1 U8830 ( .A(n23870), .B(n8222), .Y(n8229) );
  ADDFHX2 U8831 ( .A(n13371), .B(n13370), .CI(n13369), .CO(n13413), .S(n13409)
         );
  NAND2XL U8832 ( .A(n5226), .B(n9567), .Y(n5225) );
  INVXL U8833 ( .A(n5148), .Y(n5146) );
  XNOR2X1 U8834 ( .A(n4666), .B(n11971), .Y(n11965) );
  OAI21X1 U8835 ( .A0(n4410), .A1(n4092), .B0(n4090), .Y(n18353) );
  NOR2X1 U8836 ( .A(n23810), .B(n8223), .Y(n8267) );
  ADDFHX2 U8837 ( .A(n13518), .B(n13517), .CI(n13516), .CO(n13582), .S(n13544)
         );
  NAND2BXL U8838 ( .AN(n20649), .B(n6147), .Y(n20650) );
  ADDFHX2 U8839 ( .A(n16832), .B(n16831), .CI(n16830), .CO(n16837), .S(n16839)
         );
  INVXL U8840 ( .A(n9824), .Y(n5284) );
  NOR2X1 U8841 ( .A(n23858), .B(n8274), .Y(n8290) );
  NAND2X1 U8842 ( .A(n23858), .B(n8274), .Y(n8291) );
  NOR2X1 U8843 ( .A(n12784), .B(n12783), .Y(n12722) );
  OAI2BB1XL U8844 ( .A0N(n13210), .A1N(n5161), .B0(n5160), .Y(n13239) );
  NAND2XL U8845 ( .A(n13501), .B(n13502), .Y(n4494) );
  NAND2XL U8846 ( .A(n9279), .B(n4321), .Y(n4657) );
  INVXL U8847 ( .A(n9316), .Y(n5070) );
  INVXL U8848 ( .A(n4278), .Y(n4276) );
  NOR2X1 U8849 ( .A(n14925), .B(n14924), .Y(n15785) );
  NOR2X1 U8850 ( .A(n23816), .B(n8224), .Y(n8270) );
  NAND2XL U8851 ( .A(n13442), .B(n13441), .Y(n5259) );
  NAND4X1 U8852 ( .A(n25791), .B(n25789), .C(n24376), .D(n11621), .Y(n11623)
         );
  INVXL U8853 ( .A(n18361), .Y(n4410) );
  OAI21X1 U8854 ( .A0(n10301), .A1(n10496), .B0(n4358), .Y(n4357) );
  NAND2X1 U8855 ( .A(n18696), .B(n18695), .Y(n18956) );
  NAND2X1 U8856 ( .A(n4791), .B(n15017), .Y(n15042) );
  OR4XL U8857 ( .A(n23816), .B(n20374), .C(n23690), .D(n23760), .Y(n20375) );
  INVXL U8858 ( .A(n17647), .Y(n6159) );
  XOR3X2 U8859 ( .A(n17703), .B(n17704), .C(n17702), .Y(n18354) );
  INVX1 U8860 ( .A(n5865), .Y(n3169) );
  ADDFHX2 U8861 ( .A(n18596), .B(n18595), .CI(n18594), .CO(n18679), .S(n18676)
         );
  NOR2XL U8862 ( .A(n23685), .B(n7419), .Y(n7420) );
  NAND2XL U8863 ( .A(n5193), .B(n5192), .Y(n5756) );
  NAND2BXL U8864 ( .AN(n10531), .B(n5193), .Y(n5755) );
  NOR2X1 U8865 ( .A(n12786), .B(n12785), .Y(n12736) );
  NAND4X1 U8866 ( .A(n24431), .B(n24100), .C(n24355), .D(n4791), .Y(n14925) );
  NAND2X1 U8867 ( .A(n5927), .B(n5926), .Y(n17812) );
  OAI2BB1XL U8868 ( .A0N(n5540), .A1N(n10170), .B0(n5539), .Y(n10313) );
  NAND3X1 U8869 ( .A(n23816), .B(n23870), .C(n23858), .Y(n8177) );
  AOI2BB2X1 U8870 ( .B0(n10702), .B1(n10701), .A0N(n10700), .A1N(n10699), .Y(
        n25240) );
  NAND2XL U8871 ( .A(n3466), .B(n3940), .Y(n3465) );
  ADDFHX1 U8872 ( .A(n18516), .B(n18515), .CI(n18514), .CO(n18686), .S(n18683)
         );
  NAND4X1 U8873 ( .A(n23810), .B(n23844), .C(n20374), .D(n23690), .Y(n8178) );
  XOR2X1 U8874 ( .A(n5889), .B(n17796), .Y(n17859) );
  ADDFHX2 U8875 ( .A(n17818), .B(n17817), .CI(n17816), .CO(n18580), .S(n17810)
         );
  INVXL U8876 ( .A(n12215), .Y(n4016) );
  AND2X2 U8877 ( .A(n12831), .B(n12830), .Y(n12832) );
  INVX1 U8878 ( .A(n23184), .Y(n8222) );
  NAND2X1 U8879 ( .A(n24355), .B(n14969), .Y(n15012) );
  INVXL U8880 ( .A(n6668), .Y(n5554) );
  NOR2BXL U8881 ( .AN(n20652), .B(n20651), .Y(n20654) );
  OR4XL U8882 ( .A(n23870), .B(n23858), .C(n23810), .D(n23844), .Y(n20376) );
  NAND4X1 U8883 ( .A(n25129), .B(n25124), .C(n24110), .D(n18969), .Y(n18971)
         );
  NOR2X1 U8884 ( .A(n12812), .B(n12821), .Y(n12794) );
  ADDFHX1 U8885 ( .A(n13445), .B(n13444), .CI(n13443), .CO(n13489), .S(n13441)
         );
  AND2X2 U8886 ( .A(n19004), .B(n19003), .Y(n4688) );
  INVXL U8887 ( .A(n12866), .Y(n3170) );
  ADDFHX2 U8888 ( .A(n16563), .B(n16562), .CI(n16561), .CO(n16773), .S(n16768)
         );
  INVXL U8889 ( .A(n4311), .Y(n4309) );
  OAI21X2 U8890 ( .A0(n4154), .A1(n4153), .B0(n4152), .Y(n16136) );
  INVX1 U8891 ( .A(n7519), .Y(n7772) );
  OAI2BB1X1 U8892 ( .A0N(n16053), .A1N(n3635), .B0(n3631), .Y(n16059) );
  AND2XL U8893 ( .A(n14366), .B(M1_U4_U1_enc_tree_3__3__24_), .Y(n14371) );
  NOR2X1 U8894 ( .A(n18302), .B(n18301), .Y(n18305) );
  NAND2BXL U8895 ( .AN(n11920), .B(n4973), .Y(n4426) );
  INVX1 U8896 ( .A(n20169), .Y(n19309) );
  ADDFHX1 U8897 ( .A(n13719), .B(n13718), .CI(n13717), .CO(n13764), .S(n13712)
         );
  INVX1 U8898 ( .A(n7611), .Y(n7776) );
  XNOR2X1 U8899 ( .A(n21490), .B(n21489), .Y(n21496) );
  ADDFHX2 U8900 ( .A(n9333), .B(n9332), .CI(n9331), .CO(n9455), .S(n9366) );
  ADDFHX2 U8901 ( .A(n9432), .B(n9431), .CI(n9430), .CO(n9427), .S(n10086) );
  OR2X2 U8902 ( .A(n16300), .B(n16301), .Y(n5331) );
  ADDFHX2 U8903 ( .A(n7203), .B(n7202), .CI(n7201), .CO(n7266), .S(n7264) );
  AND2X2 U8904 ( .A(n17385), .B(n17384), .Y(n17386) );
  OAI21X2 U8905 ( .A0(n3813), .A1(n3812), .B0(n3811), .Y(n16194) );
  XNOR3X2 U8906 ( .A(n17004), .B(n17003), .C(n3955), .Y(n17030) );
  OAI2BB1X1 U8907 ( .A0N(n16173), .A1N(n16172), .B0(n4136), .Y(n16196) );
  OR2XL U8908 ( .A(n14187), .B(n14186), .Y(n5155) );
  INVX1 U8909 ( .A(n11789), .Y(n3900) );
  NAND2XL U8910 ( .A(n14187), .B(n14186), .Y(n5154) );
  ADDFHX2 U8911 ( .A(n7239), .B(n7238), .CI(n7237), .CO(n7262), .S(n7261) );
  ADDFHX2 U8912 ( .A(n7135), .B(n7134), .CI(n7133), .CO(n7265), .S(n7263) );
  INVXL U8913 ( .A(n5534), .Y(n5533) );
  XOR2X2 U8914 ( .A(n3794), .B(n16785), .Y(n16808) );
  NOR2X1 U8915 ( .A(n4791), .B(n15017), .Y(n15041) );
  NAND2XL U8916 ( .A(n5302), .B(n5301), .Y(n5300) );
  NAND2BXL U8917 ( .AN(n13676), .B(n13051), .Y(n5287) );
  NAND2X1 U8918 ( .A(n24050), .B(n23078), .Y(n24044) );
  ADDFHX2 U8919 ( .A(n18013), .B(n18012), .CI(n18011), .CO(n18315), .S(n18314)
         );
  INVXL U8920 ( .A(n12821), .Y(n12823) );
  NOR2XL U8921 ( .A(n5461), .B(n18134), .Y(n18216) );
  OR2XL U8922 ( .A(n10663), .B(n10662), .Y(n10665) );
  XOR2XL U8923 ( .A(n18840), .B(n17414), .Y(n17416) );
  NAND2X1 U8924 ( .A(n3419), .B(n3418), .Y(n17724) );
  OAI2BB1XL U8925 ( .A0N(n11988), .A1N(n5939), .B0(n5935), .Y(n12622) );
  NOR2X1 U8926 ( .A(n24072), .B(n19354), .Y(n19399) );
  NOR2X1 U8927 ( .A(n9163), .B(n10671), .Y(n9149) );
  NAND2BXL U8928 ( .AN(n16303), .B(n5690), .Y(n5689) );
  INVXL U8929 ( .A(n10726), .Y(n5610) );
  INVXL U8930 ( .A(n12379), .Y(n6135) );
  ADDFHX2 U8931 ( .A(n16327), .B(n16326), .CI(n16325), .CO(n17017), .S(n16300)
         );
  XNOR2X2 U8932 ( .A(n16966), .B(n4162), .Y(n17018) );
  NOR2X1 U8933 ( .A(n24390), .B(n19404), .Y(n19409) );
  XNOR3X2 U8934 ( .A(n17002), .B(n17000), .C(n17001), .Y(n3955) );
  INVXL U8935 ( .A(n18293), .Y(n5422) );
  AND2XL U8936 ( .A(M1_U4_U1_enc_tree_3__3__16_), .B(
        M1_U4_U1_enc_tree_3__3__24_), .Y(n14378) );
  NAND2X1 U8937 ( .A(n24100), .B(n14968), .Y(n14975) );
  OAI2BB1XL U8938 ( .A0N(n6509), .A1N(n6508), .B0(n5629), .Y(n6668) );
  NAND2XL U8939 ( .A(n5496), .B(n5495), .Y(n14053) );
  INVXL U8940 ( .A(n12216), .Y(n4879) );
  OAI2BB1XL U8941 ( .A0N(n14045), .A1N(n14044), .B0(n14043), .Y(n14095) );
  OR2X1 U8942 ( .A(M6_mult_x_15_n450), .B(M6_mult_x_15_n446), .Y(n10965) );
  NOR2X1 U8943 ( .A(n19308), .B(n19307), .Y(n20169) );
  AND2XL U8944 ( .A(M6_mult_x_15_n657), .B(M6_mult_x_15_n666), .Y(n10926) );
  XOR2X1 U8945 ( .A(n4871), .B(n18374), .Y(n18391) );
  NOR2X1 U8946 ( .A(n24036), .B(n22477), .Y(n24029) );
  XNOR2X1 U8947 ( .A(n5823), .B(n18588), .Y(n18579) );
  ADDFHX2 U8948 ( .A(n7212), .B(n7211), .CI(n7210), .CO(n7272), .S(n7204) );
  NAND4X1 U8949 ( .A(n25136), .B(n25132), .C(n25162), .D(n17201), .Y(n17203)
         );
  OAI21XL U8950 ( .A0(n10379), .A1(n10541), .B0(n5757), .Y(n10400) );
  NAND2XL U8951 ( .A(n6069), .B(n25862), .Y(n14231) );
  INVXL U8952 ( .A(n4974), .Y(n4973) );
  XOR3X2 U8953 ( .A(n16044), .B(n16045), .C(n16046), .Y(n16080) );
  INVX1 U8954 ( .A(n16786), .Y(n3689) );
  AND2XL U8955 ( .A(n18990), .B(n18989), .Y(n4696) );
  XNOR2X1 U8956 ( .A(n21488), .B(n21494), .Y(n21495) );
  ADDFHX2 U8957 ( .A(n7176), .B(n7175), .CI(n7174), .CO(n7205), .S(n7201) );
  NAND2XL U8958 ( .A(n6063), .B(n6061), .Y(n9511) );
  OAI2BB1XL U8959 ( .A0N(n11853), .A1N(n3914), .B0(n3912), .Y(n11839) );
  NAND2X1 U8960 ( .A(n23645), .B(n21170), .Y(n23639) );
  NAND2XL U8961 ( .A(n18698), .B(n18697), .Y(n18959) );
  NAND2X1 U8962 ( .A(n17143), .B(n17142), .Y(n17366) );
  ADDFHX2 U8963 ( .A(n7152), .B(n7151), .CI(n7150), .CO(n7202), .S(n7133) );
  ADDFHX1 U8964 ( .A(n16560), .B(n16559), .CI(n16558), .CO(n16764), .S(n16763)
         );
  NAND2XL U8965 ( .A(n4901), .B(n3448), .Y(n11869) );
  NOR2X1 U8966 ( .A(n5021), .B(n3098), .Y(n3427) );
  OR2X2 U8967 ( .A(n18698), .B(n18697), .Y(n18962) );
  NAND2BXL U8968 ( .AN(n11975), .B(n3922), .Y(n3921) );
  XNOR2X1 U8969 ( .A(n6001), .B(n12706), .Y(n12781) );
  ADDFHX1 U8970 ( .A(n11910), .B(n11909), .CI(n11908), .CO(n11935), .S(n11932)
         );
  OAI22X1 U8971 ( .A0(n8809), .A1(n3017), .B0(n3040), .B1(n8808), .Y(n8820) );
  INVXL U8972 ( .A(n5304), .Y(n5302) );
  ADDFHX2 U8973 ( .A(n9327), .B(n9326), .CI(n9325), .CO(n9392), .S(n9431) );
  INVXL U8974 ( .A(n10541), .Y(n5193) );
  ADDFHX2 U8975 ( .A(n6708), .B(n6707), .CI(n6706), .CO(n6724), .S(n6719) );
  ADDFHX2 U8976 ( .A(n6815), .B(n6814), .CI(n6813), .CO(n6905), .S(n6732) );
  ADDFHX2 U8977 ( .A(n17806), .B(n17805), .CI(n17804), .CO(n17807), .S(n17845)
         );
  NAND2XL U8978 ( .A(n17796), .B(n17797), .Y(n5926) );
  XOR3X2 U8979 ( .A(n3814), .B(n16186), .C(n16187), .Y(n16190) );
  INVXL U8980 ( .A(n6895), .Y(n5614) );
  XOR2X1 U8981 ( .A(n6894), .B(n6895), .Y(n5615) );
  NOR2X1 U8982 ( .A(n23199), .B(n23198), .Y(n10726) );
  OAI2BB1XL U8983 ( .A0N(n10533), .A1N(n10517), .B0(n10494), .Y(n10543) );
  NOR2X1 U8984 ( .A(n7721), .B(n7725), .Y(n7727) );
  NAND2BXL U8985 ( .AN(n9502), .B(n4568), .Y(n6138) );
  NAND2XL U8986 ( .A(n7576), .B(n7577), .Y(n5593) );
  ADDFHX2 U8987 ( .A(n6467), .B(n6466), .CI(n6465), .CO(n6444), .S(n6706) );
  ADDFHX2 U8988 ( .A(n6803), .B(n6802), .CI(n6801), .CO(n6893), .S(n6812) );
  NAND2X1 U8989 ( .A(n3753), .B(n3752), .Y(n17818) );
  NOR2X1 U8990 ( .A(n12792), .B(n12791), .Y(n12821) );
  NOR2X1 U8991 ( .A(n7674), .B(n7673), .Y(n7746) );
  NAND2XL U8992 ( .A(n13042), .B(n5289), .Y(n5288) );
  ADDFHX2 U8993 ( .A(n6764), .B(n6763), .CI(n6762), .CO(n6888), .S(n6809) );
  NOR2X1 U8994 ( .A(n12796), .B(n12795), .Y(n12829) );
  ADDFHX2 U8995 ( .A(n6806), .B(n6805), .CI(n6804), .CO(n6811), .S(n6813) );
  INVXL U8996 ( .A(n3913), .Y(n3912) );
  AOI2BB2XL U8997 ( .B0(n3040), .B1(n8428), .A0N(n3040), .A1N(n8475), .Y(n8542) );
  ADDFHX2 U8998 ( .A(n11991), .B(n11990), .CI(n11989), .CO(n12675), .S(n11969)
         );
  NAND2XL U8999 ( .A(n21452), .B(n21451), .Y(n21454) );
  NAND2BXL U9000 ( .AN(n9463), .B(n6062), .Y(n6061) );
  NAND2XL U9001 ( .A(n4955), .B(n4960), .Y(n4959) );
  NAND2XL U9002 ( .A(n18700), .B(n18699), .Y(n18967) );
  INVXL U9003 ( .A(n16735), .Y(n5737) );
  OR2X2 U9004 ( .A(n18700), .B(n18699), .Y(n18966) );
  NAND2XL U9005 ( .A(n11755), .B(n11754), .Y(n4901) );
  NAND2BXL U9006 ( .AN(n10402), .B(n5193), .Y(n5752) );
  AOI2BB2XL U9007 ( .B0(n3040), .B1(n8355), .A0N(n8482), .A1N(n8379), .Y(n8526) );
  ADDFHX2 U9008 ( .A(n16554), .B(n16553), .CI(n16552), .CO(n16565), .S(n16558)
         );
  ADDFHX2 U9009 ( .A(n11771), .B(n11770), .CI(n11769), .CO(n11872), .S(n11767)
         );
  XNOR2XL U9010 ( .A(n18822), .B(n18821), .Y(n18824) );
  INVXL U9011 ( .A(n18988), .Y(n18990) );
  ADDFHX2 U9012 ( .A(n6877), .B(n6876), .CI(n6875), .CO(n6891), .S(n6895) );
  AND2X1 U9013 ( .A(n19017), .B(n19016), .Y(n4697) );
  AOI2BB2XL U9014 ( .B0(n3040), .B1(n8254), .A0N(n8482), .A1N(n8327), .Y(n8536) );
  NAND2XL U9015 ( .A(n11975), .B(n3924), .Y(n3920) );
  NOR2X1 U9016 ( .A(n17396), .B(n19024), .Y(n23645) );
  AND2XL U9017 ( .A(M2_U4_U1_enc_tree_3__3__16_), .B(
        M2_U4_U1_enc_tree_3__3__24_), .Y(n10260) );
  ADDFHX2 U9018 ( .A(n17630), .B(n17629), .CI(n17628), .CO(n17850), .S(n17626)
         );
  ADDFHX2 U9019 ( .A(n16799), .B(n16798), .CI(n16797), .CO(n16828), .S(n16818)
         );
  NOR2X1 U9020 ( .A(n17135), .B(n17134), .Y(n17376) );
  INVXL U9021 ( .A(n3924), .Y(n3922) );
  NOR2X1 U9022 ( .A(n17137), .B(n17136), .Y(n17383) );
  NOR2X1 U9023 ( .A(n19025), .B(n19024), .Y(n22482) );
  AOI2BB2XL U9024 ( .B0(n3040), .B1(n8423), .A0N(n8161), .A1N(n8444), .Y(n8525) );
  NAND2BXL U9025 ( .AN(n5543), .B(n5542), .Y(n5540) );
  INVXL U9026 ( .A(n12217), .Y(n4880) );
  NAND3X1 U9027 ( .A(n24072), .B(n24390), .C(n24300), .Y(n19307) );
  INVX1 U9028 ( .A(n24401), .Y(n4792) );
  NAND2BXL U9029 ( .AN(n14014), .B(n13258), .Y(n5496) );
  NAND2BXL U9030 ( .AN(n9384), .B(n5538), .Y(n5537) );
  INVX1 U9031 ( .A(n24060), .Y(n4786) );
  NAND2X1 U9032 ( .A(n15558), .B(n14934), .Y(n14908) );
  ADDFHX2 U9033 ( .A(n16257), .B(n16256), .CI(n16255), .CO(n16265), .S(n16245)
         );
  OR2X1 U9034 ( .A(n11377), .B(n11376), .Y(n11389) );
  AOI2BB2XL U9035 ( .B0(n3040), .B1(n8235), .A0N(n8161), .A1N(n8675), .Y(n8590) );
  NAND2XL U9036 ( .A(n17952), .B(n17951), .Y(n4833) );
  ADDFHX2 U9037 ( .A(n16970), .B(n16969), .CI(n16968), .CO(n17006), .S(n17004)
         );
  NAND2X1 U9038 ( .A(n8482), .B(n8208), .Y(n8209) );
  NAND2XL U9039 ( .A(n16303), .B(n16304), .Y(n5688) );
  NAND2X1 U9040 ( .A(n8482), .B(n8200), .Y(n8201) );
  ADDFHX2 U9041 ( .A(n18382), .B(n18381), .CI(n18380), .CO(n18387), .S(n18389)
         );
  ADDFHX2 U9042 ( .A(n17667), .B(n17666), .CI(n17665), .CO(n17686), .S(n17725)
         );
  NAND2X1 U9043 ( .A(n3040), .B(n8195), .Y(n8173) );
  NAND2XL U9044 ( .A(n5936), .B(n11987), .Y(n5935) );
  OR2XL U9045 ( .A(n10679), .B(n10678), .Y(n10683) );
  NAND2X1 U9046 ( .A(n18336), .B(n18337), .Y(n3418) );
  INVX1 U9047 ( .A(n18265), .Y(n3358) );
  AOI2BB2XL U9048 ( .B0(n3040), .B1(n8237), .A0N(n3040), .A1N(n8682), .Y(n8557) );
  AOI2BB2XL U9049 ( .B0(n3040), .B1(n8297), .A0N(n8482), .A1N(n8799), .Y(n8532) );
  INVXL U9050 ( .A(n4403), .Y(n4400) );
  INVXL U9051 ( .A(n17952), .Y(n4835) );
  OR4XL U9052 ( .A(n24072), .B(n24092), .C(n24341), .D(n24295), .Y(n20135) );
  OAI22X1 U9053 ( .A0(n10368), .A1(n3831), .B0(n9345), .B1(n9780), .Y(n9365)
         );
  AOI2BB2XL U9054 ( .B0(n3040), .B1(n8307), .A0N(n3040), .A1N(n8713), .Y(n8586) );
  OR2XL U9055 ( .A(n14128), .B(n14129), .Y(n14126) );
  ADDFHX2 U9056 ( .A(n18034), .B(n18033), .CI(n18032), .CO(n18012), .S(n18096)
         );
  ADDFHX2 U9057 ( .A(n16199), .B(n16198), .CI(n16197), .CO(n16246), .S(n16195)
         );
  NAND2XL U9058 ( .A(n3867), .B(n17706), .Y(n3866) );
  INVXL U9059 ( .A(n5786), .Y(n5785) );
  INVXL U9060 ( .A(n18375), .Y(n4869) );
  OR2X2 U9061 ( .A(n6592), .B(n6591), .Y(n6556) );
  INVX1 U9062 ( .A(n14678), .Y(n14349) );
  NAND2BXL U9063 ( .AN(n18351), .B(n5877), .Y(n5876) );
  NAND2BXL U9064 ( .AN(n14250), .B(n4934), .Y(n4933) );
  INVXL U9065 ( .A(n3917), .Y(n3915) );
  NAND2BXL U9066 ( .AN(n10493), .B(n5758), .Y(n5753) );
  NAND2XL U9067 ( .A(n5810), .B(n5809), .Y(n5813) );
  NAND2XL U9068 ( .A(n5859), .B(n5545), .Y(n5857) );
  XOR2X1 U9069 ( .A(n17597), .B(n17598), .Y(n5036) );
  INVXL U9070 ( .A(n24304), .Y(n24305) );
  NAND2BXL U9071 ( .AN(n11730), .B(n4446), .Y(n4445) );
  INVXL U9072 ( .A(n24276), .Y(n4190) );
  AND2X2 U9073 ( .A(n19028), .B(n18759), .Y(n20652) );
  NOR2X1 U9074 ( .A(n18707), .B(n18706), .Y(n18988) );
  INVXL U9075 ( .A(n21450), .Y(n21452) );
  NAND2BXL U9076 ( .AN(n9501), .B(n6065), .Y(n6063) );
  NAND2X1 U9077 ( .A(n22216), .B(n23409), .Y(n22227) );
  XOR3X2 U9078 ( .A(n7178), .B(n7179), .C(n7177), .Y(n7175) );
  AND2X2 U9079 ( .A(n17399), .B(n17395), .Y(n23638) );
  ADDFHX2 U9080 ( .A(n7209), .B(n7208), .CI(n7207), .CO(n7273), .S(n7210) );
  NAND2XL U9081 ( .A(n11891), .B(n4988), .Y(n4987) );
  ADDFHX2 U9082 ( .A(n7279), .B(n7278), .CI(n7277), .CO(n7454), .S(n7271) );
  ADDFHX2 U9083 ( .A(n7518), .B(n7517), .CI(n7516), .CO(n7608), .S(n7492) );
  ADDFHX2 U9084 ( .A(n7598), .B(n7597), .CI(n7596), .CO(n7606), .S(n7609) );
  OAI21XL U9085 ( .A0(n5444), .A1(n5442), .B0(n5440), .Y(n18510) );
  ADDFHX2 U9086 ( .A(n18587), .B(n18586), .CI(n18585), .CO(n18594), .S(n18592)
         );
  NAND2XL U9087 ( .A(n5517), .B(n6065), .Y(n6064) );
  NOR2X1 U9088 ( .A(n7717), .B(n7716), .Y(n7725) );
  NOR2X1 U9089 ( .A(n7740), .B(n7739), .Y(n7791) );
  NAND2X1 U9090 ( .A(n7740), .B(n7739), .Y(n7790) );
  INVX1 U9091 ( .A(n7816), .Y(n7817) );
  INVXL U9092 ( .A(n11693), .Y(n4960) );
  NAND2XL U9093 ( .A(n5619), .B(n6531), .Y(n5618) );
  INVXL U9094 ( .A(n3764), .Y(n3763) );
  ADDFHX2 U9095 ( .A(n6702), .B(n6701), .CI(n6700), .CO(n6707), .S(n6709) );
  OAI2BB1XL U9096 ( .A0N(n5323), .A1N(n5962), .B0(n4751), .Y(n5322) );
  INVXL U9097 ( .A(n13600), .Y(n5289) );
  ADDFHX1 U9098 ( .A(n6448), .B(n6447), .CI(n6446), .CO(n6440), .S(n6708) );
  NAND2BXL U9099 ( .AN(n9223), .B(n6065), .Y(n6060) );
  XOR3X2 U9100 ( .A(n6770), .B(n6769), .C(n6768), .Y(n6815) );
  OAI21XL U9101 ( .A0(n6769), .A1(n6770), .B0(n6768), .Y(n3498) );
  ADDFHX2 U9102 ( .A(n6800), .B(n6799), .CI(n6798), .CO(n6801), .S(n6805) );
  NAND2XL U9103 ( .A(n11717), .B(n11716), .Y(n3644) );
  OAI22X1 U9104 ( .A0(n19938), .A1(n3100), .B0(n3041), .B1(n19937), .Y(n19949)
         );
  NAND2BXL U9105 ( .AN(n10402), .B(n5758), .Y(n5757) );
  NAND2BXL U9106 ( .AN(n11875), .B(n5974), .Y(n5973) );
  ADDFHX2 U9107 ( .A(n7126), .B(n7125), .CI(n7124), .CO(n7248), .S(n7244) );
  ADDFHX2 U9108 ( .A(n7104), .B(n7103), .CI(n7102), .CO(n7151), .S(n7123) );
  NAND2XL U9109 ( .A(n16099), .B(n4780), .Y(n6150) );
  NAND2XL U9110 ( .A(n17632), .B(n3823), .Y(n3821) );
  NAND2BXL U9111 ( .AN(n10531), .B(n5758), .Y(n5754) );
  INVXL U9112 ( .A(n12177), .Y(n6004) );
  OAI21XL U9113 ( .A0(n16960), .A1(n5329), .B0(n5328), .Y(n16324) );
  OAI21XL U9114 ( .A0(n16960), .A1(n5947), .B0(n5946), .Y(n16986) );
  OAI2BB1XL U9115 ( .A0N(n17568), .A1N(n3406), .B0(n3402), .Y(n17615) );
  NAND2XL U9116 ( .A(n18076), .B(n18077), .Y(n6126) );
  OAI22XL U9117 ( .A0(n14076), .A1(n14227), .B0(n14249), .B1(n4298), .Y(n14096) );
  OAI2BB1XL U9118 ( .A0N(n10496), .A1N(n9504), .B0(n4808), .Y(n10509) );
  XOR2X1 U9119 ( .A(n11854), .B(n3917), .Y(n3916) );
  INVXL U9120 ( .A(n3635), .Y(n3633) );
  ADDFHX2 U9121 ( .A(n16993), .B(n16992), .CI(n16991), .CO(n17022), .S(n17024)
         );
  NAND2BXL U9122 ( .AN(n11988), .B(n5937), .Y(n5936) );
  XOR2X1 U9123 ( .A(n16052), .B(n3635), .Y(n3634) );
  OR2XL U9124 ( .A(n10692), .B(n10676), .Y(n9188) );
  NAND2BXL U9125 ( .AN(n11977), .B(n5371), .Y(n5370) );
  NAND2BXL U9126 ( .AN(n9960), .B(n9904), .Y(n9905) );
  OR2X2 U9127 ( .A(n9906), .B(n9904), .Y(n4312) );
  INVX2 U9128 ( .A(n14121), .Y(n13258) );
  AND2XL U9129 ( .A(n18199), .B(n18198), .Y(n18203) );
  NAND2XL U9130 ( .A(n4420), .B(n11846), .Y(n4419) );
  INVXL U9131 ( .A(n12445), .Y(n11815) );
  XNOR3X2 U9132 ( .A(n17972), .B(n17971), .C(n3410), .Y(n4403) );
  ADDFHX2 U9133 ( .A(n17991), .B(n17990), .CI(n17989), .CO(n17983), .S(n18013)
         );
  OAI21XL U9134 ( .A0(n17971), .A1(n17972), .B0(n3410), .Y(n5816) );
  XNOR2X1 U9135 ( .A(n3751), .B(n17773), .Y(n17809) );
  XOR3X2 U9136 ( .A(n16119), .B(n16118), .C(n16120), .Y(n16150) );
  XOR2X1 U9137 ( .A(n16172), .B(n16173), .Y(n3370) );
  NAND2XL U9138 ( .A(n6080), .B(n4087), .Y(n6077) );
  OAI2BB1X2 U9139 ( .A0N(n5804), .A1N(n16427), .B0(n5803), .Y(n16798) );
  NAND2BXL U9140 ( .AN(n6080), .B(n4171), .Y(n6079) );
  ADDFHX2 U9141 ( .A(n15992), .B(n15991), .CI(n15990), .CO(n16043), .S(n15993)
         );
  NAND2XL U9142 ( .A(n16160), .B(n16159), .Y(n5954) );
  NOR2X1 U9143 ( .A(n11576), .B(n13006), .Y(n13003) );
  AND2X2 U9144 ( .A(n13006), .B(n11576), .Y(n24043) );
  XOR2X1 U9145 ( .A(n12107), .B(n3846), .Y(n3381) );
  OAI21XL U9146 ( .A0(n6076), .A1(n9892), .B0(n4335), .Y(n4332) );
  NAND2XL U9147 ( .A(n5725), .B(n16967), .Y(n5722) );
  NAND2X2 U9148 ( .A(n4667), .B(n14120), .Y(n14121) );
  NAND2BXL U9149 ( .AN(n13792), .B(n13203), .Y(n5503) );
  XOR2X1 U9150 ( .A(n6983), .B(n6984), .Y(n4553) );
  INVXL U9151 ( .A(n12185), .Y(n3993) );
  XOR2X1 U9152 ( .A(n11976), .B(n5373), .Y(n5372) );
  INVXL U9153 ( .A(n12583), .Y(n4046) );
  NAND2BXL U9154 ( .AN(n9383), .B(n5536), .Y(n5535) );
  INVXL U9155 ( .A(n17067), .Y(n5095) );
  NAND2XL U9156 ( .A(n5884), .B(n17739), .Y(n5883) );
  NAND2BXL U9157 ( .AN(n6532), .B(n5575), .Y(n5619) );
  NAND2XL U9158 ( .A(n18281), .B(n18282), .Y(n5423) );
  NAND2BXL U9159 ( .AN(n16974), .B(n4097), .Y(n4096) );
  INVXL U9160 ( .A(n18352), .Y(n5877) );
  OAI21X1 U9161 ( .A0(n15955), .A1(n16960), .B0(n3618), .Y(n15992) );
  NAND2BXL U9162 ( .AN(n17940), .B(n4392), .Y(n4391) );
  NAND2XL U9163 ( .A(n18351), .B(n18352), .Y(n5875) );
  NOR2X1 U9164 ( .A(n9128), .B(n9127), .Y(n10671) );
  NAND2X1 U9165 ( .A(n11580), .B(n13007), .Y(n11576) );
  INVXL U9166 ( .A(n3870), .Y(n3867) );
  INVXL U9167 ( .A(n17972), .Y(n5818) );
  AND2XL U9168 ( .A(M3_U3_U1_enc_tree_3__3__16_), .B(
        M3_U3_U1_enc_tree_3__3__24_), .Y(n12955) );
  XNOR2X1 U9169 ( .A(n4393), .B(n4031), .Y(n3410) );
  OR2XL U9170 ( .A(n6590), .B(n6589), .Y(n6562) );
  NAND2BXL U9171 ( .AN(n14058), .B(n13203), .Y(n5495) );
  NAND2X1 U9172 ( .A(n3018), .B(n3685), .Y(n3684) );
  ADDFHX1 U9173 ( .A(n18254), .B(n18253), .CI(n18252), .CO(n18287), .S(n18255)
         );
  NOR2X1 U9174 ( .A(n9113), .B(n9112), .Y(n10680) );
  NAND2XL U9175 ( .A(n17919), .B(n5811), .Y(n5812) );
  INVXL U9176 ( .A(n17919), .Y(n5810) );
  NAND2XL U9177 ( .A(n4912), .B(n12643), .Y(n4911) );
  NOR2X1 U9178 ( .A(n9135), .B(n9134), .Y(n10677) );
  NAND2XL U9179 ( .A(n17720), .B(n3765), .Y(n3762) );
  INVXL U9180 ( .A(n6698), .Y(n5625) );
  NAND2BXL U9181 ( .AN(n9960), .B(n10494), .Y(n9442) );
  NOR2X1 U9182 ( .A(n21404), .B(n21403), .Y(n22216) );
  AOI2BB2XL U9183 ( .B0(n15008), .B1(n15175), .A0N(n15190), .A1N(n15207), .Y(
        n15296) );
  NAND4X1 U9184 ( .A(n21441), .B(n21440), .C(n21439), .D(n21438), .Y(n21442)
         );
  OR2XL U9185 ( .A(n11798), .B(n5789), .Y(n5787) );
  AND2XL U9186 ( .A(n11798), .B(n5789), .Y(n5786) );
  NAND2XL U9187 ( .A(n11922), .B(n3660), .Y(n3659) );
  INVXL U9188 ( .A(n11922), .Y(n3662) );
  NAND2BXL U9189 ( .AN(n9960), .B(n25885), .Y(n9324) );
  NAND2XL U9190 ( .A(n7140), .B(n7141), .Y(n5563) );
  XNOR2X1 U9191 ( .A(n10324), .B(n9901), .Y(n9774) );
  NOR2XL U9192 ( .A(n10324), .B(n9841), .Y(M2_U3_U1_or2_tree_0__1__20_) );
  NAND2BXL U9193 ( .AN(n17534), .B(n5863), .Y(n5862) );
  INVXL U9194 ( .A(n5782), .Y(n5777) );
  OR2XL U9195 ( .A(n23413), .B(n21493), .Y(n21492) );
  NOR2X1 U9196 ( .A(n23394), .B(n21486), .Y(n21491) );
  INVXL U9197 ( .A(n4423), .Y(n4420) );
  XOR2X1 U9198 ( .A(n11835), .B(n4925), .Y(n12442) );
  XOR3X2 U9199 ( .A(n4423), .B(n4422), .C(n11845), .Y(n12437) );
  XOR2X1 U9200 ( .A(n10494), .B(M2_U4_U1_or2_inv_0__22_), .Y(n9362) );
  NAND2XL U9201 ( .A(n3403), .B(n17567), .Y(n3402) );
  OAI2BB1XL U9202 ( .A0N(n17775), .A1N(n4883), .B0(n4650), .Y(n17821) );
  NAND2X1 U9203 ( .A(n23402), .B(n21445), .Y(n21480) );
  NAND2X1 U9204 ( .A(n14362), .B(n14361), .Y(n4677) );
  INVXL U9205 ( .A(n11874), .Y(n5974) );
  NAND2XL U9206 ( .A(n11875), .B(n11874), .Y(n5972) );
  NAND2XL U9207 ( .A(n12697), .B(n5994), .Y(n5993) );
  NOR2X1 U9208 ( .A(n18711), .B(n18710), .Y(n19015) );
  NAND2X1 U9209 ( .A(n17179), .B(n17400), .Y(n17395) );
  AND2X2 U9210 ( .A(n18726), .B(n18725), .Y(n4699) );
  ADDFHX1 U9211 ( .A(n11913), .B(n4774), .CI(n11911), .CO(n11961), .S(n11909)
         );
  INVXL U9212 ( .A(n4990), .Y(n4988) );
  OAI22XL U9213 ( .A0(n10660), .A1(n9874), .B0(n10659), .B1(n9863), .Y(n9346)
         );
  NOR2X1 U9214 ( .A(n7387), .B(n7848), .Y(n7869) );
  NAND2X1 U9215 ( .A(n7387), .B(n7848), .Y(n7836) );
  INVXL U9216 ( .A(n10362), .Y(n5192) );
  ADDFHX1 U9217 ( .A(n11685), .B(n11684), .CI(n11683), .CO(n11711), .S(n11737)
         );
  INVXL U9218 ( .A(n11686), .Y(n5323) );
  OAI21XL U9219 ( .A0(n18550), .A1(n5441), .B0(n18549), .Y(n5440) );
  INVXL U9220 ( .A(n18550), .Y(n5442) );
  ADDFHX2 U9221 ( .A(n7583), .B(n7582), .CI(n7581), .CO(n7652), .S(n7575) );
  NAND2X1 U9222 ( .A(n3041), .B(n19314), .Y(n19293) );
  INVXL U9223 ( .A(n16820), .Y(n3779) );
  NAND2X1 U9224 ( .A(n19564), .B(n19333), .Y(n19300) );
  NAND2XL U9225 ( .A(n17771), .B(n4373), .Y(n4370) );
  OR2XL U9226 ( .A(n4373), .B(n17771), .Y(n4371) );
  XOR2X1 U9227 ( .A(n3417), .B(n5782), .Y(n5781) );
  INVX1 U9228 ( .A(n16449), .Y(n4113) );
  INVXL U9229 ( .A(n18557), .Y(n4247) );
  AND2XL U9230 ( .A(n12169), .B(n5509), .Y(n12166) );
  XOR2X1 U9231 ( .A(n3643), .B(n3642), .Y(n11889) );
  NOR2XL U9232 ( .A(n17607), .B(n4409), .Y(n4489) );
  AND2X2 U9233 ( .A(n6344), .B(n6343), .Y(n6760) );
  NAND2XL U9234 ( .A(n18724), .B(n18723), .Y(n18725) );
  NAND2BXL U9235 ( .AN(n16382), .B(n3179), .Y(n3616) );
  INVXL U9236 ( .A(n9906), .Y(n5536) );
  NOR2BXL U9237 ( .AN(n5512), .B(n25862), .Y(M1_U4_U1_or2_tree_0__1__16_) );
  NAND2BXL U9238 ( .AN(n11851), .B(n3383), .Y(n3918) );
  XOR2X2 U9239 ( .A(n14156), .B(n4502), .Y(n4503) );
  INVXL U9240 ( .A(n10387), .Y(n10365) );
  INVXL U9241 ( .A(n4171), .Y(n4087) );
  AND2XL U9242 ( .A(n17268), .B(M5_U3_U1_enc_tree_3__3__24_), .Y(n17272) );
  NOR2X1 U9243 ( .A(n7391), .B(n7849), .Y(n7387) );
  NAND2XL U9244 ( .A(n17534), .B(n5864), .Y(n5861) );
  INVXL U9245 ( .A(n5864), .Y(n5863) );
  AND2XL U9246 ( .A(n18798), .B(M4_U3_U1_enc_tree_3__3__24_), .Y(n18803) );
  INVXL U9247 ( .A(n5909), .Y(n5906) );
  NAND2BXL U9248 ( .AN(n17568), .B(n3404), .Y(n3403) );
  NAND2XL U9249 ( .A(n5066), .B(n5064), .Y(n5063) );
  XOR2X1 U9250 ( .A(n17567), .B(n3405), .Y(n17572) );
  INVX1 U9251 ( .A(n12357), .Y(n3383) );
  INVXL U9252 ( .A(n4926), .Y(n4924) );
  INVXL U9253 ( .A(n5797), .Y(n5794) );
  NAND2XL U9254 ( .A(n3179), .B(n3623), .Y(n3622) );
  AND2XL U9255 ( .A(M2_U4_U1_or2_inv_0__18_), .B(n10337), .Y(n5742) );
  NAND2BXL U9256 ( .AN(n17730), .B(n5797), .Y(n5795) );
  INVXL U9257 ( .A(n5672), .Y(n5670) );
  NOR2X1 U9258 ( .A(n18761), .B(n19031), .Y(n18760) );
  XOR2X2 U9259 ( .A(M2_a_18_), .B(n5202), .Y(n9215) );
  NAND2BXL U9260 ( .AN(n11666), .B(n3732), .Y(n3731) );
  INVXL U9261 ( .A(n4075), .Y(n4074) );
  INVXL U9262 ( .A(n5444), .Y(n5441) );
  INVXL U9263 ( .A(n9892), .Y(n4333) );
  OAI21X1 U9264 ( .A0(n15997), .A1(n5835), .B0(n3701), .Y(n16055) );
  INVXL U9265 ( .A(n6699), .Y(n5626) );
  NAND2X1 U9266 ( .A(n5325), .B(n5324), .Y(n11686) );
  NOR2BXL U9267 ( .AN(n5512), .B(M1_b_12_), .Y(M1_U4_U1_enc_tree_1__1__18_) );
  NAND2XL U9268 ( .A(n5894), .B(n18453), .Y(n18469) );
  XNOR2X1 U9269 ( .A(n14266), .B(n14228), .Y(n4298) );
  OAI2BB1XL U9270 ( .A0N(n12760), .A1N(n12759), .B0(n12758), .Y(n12801) );
  NAND2BXL U9271 ( .AN(n16869), .B(n5945), .Y(n5944) );
  OAI21XL U9272 ( .A0(n12617), .A1(n12616), .B0(n3964), .Y(n12614) );
  INVXL U9273 ( .A(n17706), .Y(n3869) );
  INVXL U9274 ( .A(n4099), .Y(n4097) );
  INVXL U9275 ( .A(n4394), .Y(n4392) );
  NOR2X1 U9276 ( .A(n11584), .B(n13009), .Y(n11580) );
  NAND2XL U9277 ( .A(n11666), .B(n3734), .Y(n3730) );
  NOR2X1 U9278 ( .A(n17180), .B(n17402), .Y(n17179) );
  ADDFHX2 U9279 ( .A(n7230), .B(n7229), .CI(n7228), .CO(n7275), .S(n7208) );
  INVXL U9280 ( .A(n3697), .Y(n3695) );
  NOR2X1 U9281 ( .A(n14433), .B(n14707), .Y(n14693) );
  NAND2XL U9282 ( .A(n4438), .B(n4437), .Y(n4436) );
  INVX2 U9283 ( .A(n5725), .Y(n3176) );
  ADDFHX2 U9284 ( .A(n6797), .B(n6796), .CI(n6795), .CO(n6802), .S(n6768) );
  INVXL U9285 ( .A(n5811), .Y(n5809) );
  NAND2BXL U9286 ( .AN(n16103), .B(n3179), .Y(n3620) );
  NAND4X1 U9287 ( .A(n9138), .B(n9137), .C(n9136), .D(n25210), .Y(n10681) );
  XOR2X1 U9288 ( .A(n4751), .B(n5964), .Y(n5963) );
  NAND3X1 U9289 ( .A(n9144), .B(n9143), .C(n14432), .Y(n10686) );
  NAND2BXL U9290 ( .AN(n12644), .B(n4914), .Y(n4912) );
  NAND2BXL U9291 ( .AN(n16497), .B(n5847), .Y(n5846) );
  INVXL U9292 ( .A(n4440), .Y(n4438) );
  NOR2X2 U9293 ( .A(n5910), .B(n4847), .Y(n5909) );
  NAND2BXL U9294 ( .AN(n11793), .B(n4134), .Y(n4135) );
  INVX8 U9295 ( .A(n4288), .Y(n14228) );
  NAND2BXL U9296 ( .AN(n18041), .B(n5458), .Y(n5457) );
  INVXL U9297 ( .A(n17591), .Y(n5873) );
  INVXL U9298 ( .A(n4041), .Y(n4039) );
  INVXL U9299 ( .A(n16967), .Y(n5724) );
  INVXL U9300 ( .A(n17607), .Y(n4487) );
  INVXL U9301 ( .A(n4488), .Y(n4409) );
  BUFX3 U9302 ( .A(n23222), .Y(M2_mult_x_15_n1669) );
  INVXL U9303 ( .A(n6104), .Y(n6101) );
  XOR2X1 U9304 ( .A(n3969), .B(n3968), .Y(n12694) );
  NAND2XL U9305 ( .A(n4909), .B(n4908), .Y(n4907) );
  INVXL U9306 ( .A(n3875), .Y(n3873) );
  NAND2XL U9307 ( .A(n3965), .B(n5941), .Y(n5940) );
  NAND2XL U9308 ( .A(n6104), .B(n6103), .Y(n6102) );
  AND2XL U9309 ( .A(M5_U3_U1_enc_tree_3__3__16_), .B(
        M5_U3_U1_enc_tree_3__3__24_), .Y(n17278) );
  NAND2BXL U9310 ( .AN(n17903), .B(n3104), .Y(n5819) );
  INVXL U9311 ( .A(n16960), .Y(n5945) );
  NOR4XL U9312 ( .A(n23822), .B(n23865), .C(n23782), .D(n23862), .Y(n7418) );
  BUFX8 U9313 ( .A(n10659), .Y(n3178) );
  AND2XL U9314 ( .A(M0_U4_U1_enc_tree_3__3__16_), .B(
        M0_U4_U1_enc_tree_3__3__24_), .Y(n7341) );
  INVX1 U9315 ( .A(M2_a_22_), .Y(n9221) );
  AND2XL U9316 ( .A(n7330), .B(M0_U3_U1_enc_tree_3__3__24_), .Y(n7334) );
  NAND2XL U9317 ( .A(n5941), .B(n4997), .Y(n4996) );
  XOR2X1 U9318 ( .A(M1_b_18_), .B(M1_b_19_), .Y(n13427) );
  NAND2BXL U9319 ( .AN(n18433), .B(n5896), .Y(n5895) );
  NAND2XL U9320 ( .A(n5463), .B(n18500), .Y(n18435) );
  NAND2BXL U9321 ( .AN(n11721), .B(n5326), .Y(n5325) );
  NAND2X1 U9322 ( .A(n11588), .B(n13010), .Y(n11584) );
  NAND2BXL U9323 ( .AN(n17966), .B(n3855), .Y(n3854) );
  NAND2XL U9324 ( .A(n5732), .B(n5760), .Y(n5759) );
  NAND2X1 U9325 ( .A(n14437), .B(n14704), .Y(n14433) );
  CLKINVX3 U9326 ( .A(M2_a_12_), .Y(n5250) );
  OAI2BB1XL U9327 ( .A0N(n12746), .A1N(n12715), .B0(n12732), .Y(n12753) );
  NAND4X1 U9328 ( .A(n14456), .B(n14432), .C(n14431), .D(n14430), .Y(n14716)
         );
  NOR2BXL U9329 ( .AN(M2_U4_U1_or2_inv_0__26_), .B(M2_b_4_), .Y(
        M2_U4_U1_enc_tree_1__1__26_) );
  OAI21XL U9330 ( .A0(n3046), .A1(n3542), .B0(n3540), .Y(n7099) );
  INVXL U9331 ( .A(n3734), .Y(n3732) );
  NAND3X1 U9332 ( .A(n14405), .B(n14404), .C(n14403), .Y(n14715) );
  NOR2BXL U9333 ( .AN(M2_U4_U1_or2_inv_0__26_), .B(M2_b_7_), .Y(
        M2_U4_U1_or2_tree_0__1__24_) );
  INVXL U9334 ( .A(n5887), .Y(n5885) );
  INVX1 U9335 ( .A(M1_b_2_), .Y(n5168) );
  NAND2XL U9336 ( .A(n11750), .B(n11751), .Y(n3652) );
  NAND2XL U9337 ( .A(n5734), .B(n4165), .Y(n5733) );
  INVXL U9338 ( .A(n15976), .Y(n6121) );
  NAND2BXL U9339 ( .AN(n11722), .B(n5415), .Y(n5790) );
  NAND2XL U9340 ( .A(n5732), .B(n5734), .Y(n5731) );
  NAND2X1 U9341 ( .A(n7393), .B(n7847), .Y(n7391) );
  NAND2XL U9342 ( .A(n3904), .B(n12519), .Y(n12562) );
  AND2XL U9343 ( .A(M1_U3_U1_enc_tree_3__3__16_), .B(
        M1_U3_U1_enc_tree_3__3__24_), .Y(n14379) );
  NAND2BXL U9344 ( .AN(n12618), .B(n3965), .Y(n3964) );
  INVXL U9345 ( .A(n11781), .Y(n4991) );
  CMPR22X1 U9346 ( .A(n11676), .B(n11675), .CO(n11725), .S(n11731) );
  INVXL U9347 ( .A(n24348), .Y(n6131) );
  XOR2X1 U9348 ( .A(n17993), .B(n3440), .Y(n18021) );
  INVXL U9349 ( .A(n20788), .Y(n3771) );
  INVXL U9350 ( .A(n12206), .Y(n4739) );
  NAND2X1 U9351 ( .A(n17181), .B(n17403), .Y(n17180) );
  OAI22XL U9352 ( .A0(n12065), .A1(n12598), .B0(n12342), .B1(n12030), .Y(
        n12078) );
  NAND2BXL U9353 ( .AN(n7052), .B(n5122), .Y(n5113) );
  NAND2X1 U9354 ( .A(n9064), .B(n13507), .Y(n23222) );
  NAND2XL U9355 ( .A(n6013), .B(n16965), .Y(n6011) );
  CLKINVX4 U9356 ( .A(M1_b_0_), .Y(n3181) );
  NOR2XL U9357 ( .A(n25884), .B(n4431), .Y(M3_U3_U1_enc_tree_1__1__16_) );
  NAND2XL U9358 ( .A(n5675), .B(n5674), .Y(n5673) );
  NAND2BXL U9359 ( .AN(n6824), .B(n5122), .Y(n5121) );
  BUFX8 U9360 ( .A(n9058), .Y(M2_mult_x_15_a_1_) );
  AOI2BB2XL U9361 ( .B0(n23116), .B1(n21790), .A0N(n21628), .A1N(n21791), .Y(
        n21691) );
  OR2XL U9362 ( .A(M4_U4_U1_enc_tree_2__2__16_), .B(
        M4_U4_U1_enc_tree_2__2__24_), .Y(n26146) );
  OAI21X2 U9363 ( .A0(n12340), .A1(n3728), .B0(n3727), .Y(n11750) );
  OAI21XL U9364 ( .A0(n18659), .A1(n4200), .B0(n4199), .Y(n18634) );
  ADDFHX1 U9365 ( .A(n3110), .B(n11646), .CI(n11645), .CO(n11660), .S(n11724)
         );
  OAI2BB1XL U9366 ( .A0N(n12222), .A1N(n12352), .B0(n12233), .Y(n11987) );
  OAI21XL U9367 ( .A0(n16341), .A1(n16686), .B0(n3936), .Y(n16355) );
  OAI2BB1XL U9368 ( .A0N(n12616), .A1N(n12618), .B0(n25884), .Y(n12697) );
  NAND2XL U9369 ( .A(n12635), .B(n12633), .Y(n3904) );
  NAND2BXL U9370 ( .AN(n6977), .B(n5122), .Y(n5112) );
  NAND3X1 U9371 ( .A(n9044), .B(n5763), .C(n5762), .Y(M2_a_14_) );
  XOR2X1 U9372 ( .A(n5960), .B(n16289), .Y(n4126) );
  NOR2BX2 U9373 ( .AN(n9054), .B(n3264), .Y(n3263) );
  NOR2BX2 U9374 ( .AN(n9078), .B(n4322), .Y(M2_U4_U1_or2_inv_0__22_) );
  NOR2X1 U9375 ( .A(n18763), .B(n19034), .Y(n18762) );
  NOR2X1 U9376 ( .A(n14441), .B(n14705), .Y(n14437) );
  INVXL U9377 ( .A(n12525), .Y(n4909) );
  ADDFHX1 U9378 ( .A(n6333), .B(n6332), .CI(n6331), .CO(n6357), .S(n6353) );
  NAND2BXL U9379 ( .AN(n7546), .B(n5122), .Y(n5108) );
  NOR2X1 U9380 ( .A(n11592), .B(n13012), .Y(n11588) );
  NAND2XL U9381 ( .A(n11881), .B(n3114), .Y(n3640) );
  OR2XL U9382 ( .A(M3_U4_U1_or2_tree_1__2__16_), .B(
        M3_U4_U1_or2_tree_1__2__24_), .Y(n26155) );
  INVXL U9383 ( .A(n3857), .Y(n3855) );
  NAND2XL U9384 ( .A(n17966), .B(n3857), .Y(n3853) );
  OAI2BB1XL U9385 ( .A0N(n6613), .A1N(n6608), .B0(n25867), .Y(n7233) );
  NAND2BXL U9386 ( .AN(n7292), .B(n5122), .Y(n5118) );
  INVXL U9387 ( .A(n24239), .Y(n3974) );
  OAI21X1 U9388 ( .A0(n7190), .A1(n7288), .B0(n3577), .Y(n7192) );
  NAND4BX2 U9389 ( .AN(n25150), .B(n5253), .C(n5252), .D(n5251), .Y(M2_a_12_)
         );
  OAI22X1 U9390 ( .A0(n11654), .A1(n12598), .B0(n12342), .B1(n3738), .Y(n11774) );
  NOR2X1 U9391 ( .A(n7395), .B(n7845), .Y(n7393) );
  OAI21X1 U9392 ( .A0(n4169), .A1(n16686), .B0(n4168), .Y(n16071) );
  INVXL U9393 ( .A(n4908), .Y(n4906) );
  NAND3X1 U9394 ( .A(n9141), .B(n9140), .C(n14405), .Y(n10684) );
  INVX4 U9395 ( .A(n6076), .Y(n3182) );
  NAND2XL U9396 ( .A(n25870), .B(n5110), .Y(n7714) );
  NOR2X1 U9397 ( .A(n13002), .B(n13001), .Y(n19024) );
  NOR2X1 U9398 ( .A(n17182), .B(n17405), .Y(n17181) );
  NAND2XL U9399 ( .A(n3451), .B(n5122), .Y(n5106) );
  NAND2XL U9400 ( .A(n3424), .B(n3637), .Y(n3619) );
  NAND2BXL U9401 ( .AN(n7563), .B(n5122), .Y(n5107) );
  INVXL U9402 ( .A(n12632), .Y(n4915) );
  NAND2BXL U9403 ( .AN(n7089), .B(n5122), .Y(n5119) );
  ADDFX2 U9404 ( .A(M4_mult_x_15_n1680), .B(n3190), .CI(n18427), .CO(n18442), 
        .S(n18495) );
  OAI22X1 U9405 ( .A0(n17060), .A1(n16102), .B0(n17061), .B1(n16087), .Y(
        n16106) );
  INVXL U9406 ( .A(n12635), .Y(n4916) );
  AND2XL U9407 ( .A(M0_U3_U1_enc_tree_3__3__16_), .B(
        M0_U3_U1_enc_tree_3__3__24_), .Y(n7342) );
  INVXL U9408 ( .A(n6008), .Y(n4504) );
  INVXL U9409 ( .A(n5893), .Y(n5896) );
  NAND2X1 U9410 ( .A(n11536), .B(learning_rate[12]), .Y(n4273) );
  OR2XL U9411 ( .A(n25870), .B(n6299), .Y(M0_U3_U1_or2_tree_0__1__12_) );
  OAI2BB1XL U9412 ( .A0N(n17061), .A1N(n17060), .B0(n17039), .Y(n17068) );
  NOR2XL U9413 ( .A(n25864), .B(M1_a_19_), .Y(M1_U3_U1_enc_tree_1__1__12_) );
  NAND2X1 U9414 ( .A(n8113), .B(n8156), .Y(n8159) );
  AND2XL U9415 ( .A(n7829), .B(n7828), .Y(n7830) );
  AOI21XL U9416 ( .A0(n4002), .A1(n3740), .B0(n3639), .Y(
        M3_U3_U1_enc_tree_0__1__26_) );
  INVXL U9417 ( .A(n4777), .Y(M3_a_2_) );
  NAND2BX1 U9418 ( .AN(n7166), .B(n3578), .Y(n3577) );
  NAND2XL U9419 ( .A(M4_a_0_), .B(n6035), .Y(n6034) );
  NAND2XL U9420 ( .A(n20743), .B(n25206), .Y(n4849) );
  NAND2X2 U9421 ( .A(n3796), .B(n15949), .Y(n16867) );
  NOR2XL U9422 ( .A(M3_mult_x_15_b_9_), .B(n5430), .Y(
        M4_U4_U1_enc_tree_1__1__22_) );
  AND2XL U9423 ( .A(n3110), .B(n3637), .Y(n16495) );
  NAND2BXL U9424 ( .AN(n3110), .B(n12519), .Y(n12132) );
  AND2XL U9425 ( .A(M4_U4_U1_enc_tree_1__1__12_), .B(
        M4_U4_U1_enc_tree_1__1__14_), .Y(n25893) );
  INVXL U9426 ( .A(n16938), .Y(n5675) );
  INVXL U9427 ( .A(n5729), .Y(n4164) );
  INVXL U9428 ( .A(n5061), .Y(n5060) );
  BUFX8 U9429 ( .A(n17099), .Y(n16317) );
  INVXL U9430 ( .A(n13695), .Y(n6055) );
  INVXL U9431 ( .A(n3937), .Y(n3935) );
  INVXL U9432 ( .A(n12119), .Y(n3874) );
  INVXL U9433 ( .A(n4876), .Y(n5898) );
  NOR2X1 U9434 ( .A(n9087), .B(n25907), .Y(n3264) );
  INVXL U9435 ( .A(n12519), .Y(n4513) );
  OAI2BB1XL U9436 ( .A0N(n18653), .A1N(n18652), .B0(n18638), .Y(n18661) );
  NAND2XL U9437 ( .A(n5705), .B(n6124), .Y(n6123) );
  NAND2XL U9438 ( .A(n20937), .B(n4772), .Y(n4851) );
  INVXL U9439 ( .A(n12542), .Y(n4437) );
  INVX1 U9440 ( .A(n12105), .Y(n3382) );
  AND2XL U9441 ( .A(n23080), .B(n23079), .Y(n23083) );
  INVXL U9442 ( .A(n16965), .Y(n4166) );
  NOR2XL U9443 ( .A(n12732), .B(n4918), .Y(M3_U3_U1_enc_tree_1__1__12_) );
  INVXL U9444 ( .A(n16943), .Y(n4165) );
  NOR2X1 U9445 ( .A(n18755), .B(n18754), .Y(n19031) );
  OAI21XL U9446 ( .A0(n17512), .A1(n2978), .B0(n18721), .Y(n17540) );
  NOR2XL U9447 ( .A(n11485), .B(n3740), .Y(M3_U3_U1_enc_tree_1__1__24_) );
  NAND2XL U9448 ( .A(n20734), .B(n3111), .Y(n5337) );
  AOI22XL U9449 ( .A0(n25754), .A1(sigma11[3]), .B0(sigma12[3]), .B1(n20748), 
        .Y(n20749) );
  AOI21XL U9450 ( .A0(n4431), .A1(M3_U3_U1_or2_inv_0__18_), .B0(n5045), .Y(
        M3_U3_U1_enc_tree_0__1__18_) );
  AOI22XL U9451 ( .A0(n25763), .A1(n25932), .B0(n25754), .B1(n26445), .Y(
        n20339) );
  NOR2XL U9452 ( .A(n12265), .B(n3639), .Y(M3_U3_U1_enc_tree_1__1__26_) );
  AOI22XL U9453 ( .A0(n25763), .A1(n26031), .B0(n25754), .B1(n26444), .Y(
        n24134) );
  AOI22XL U9454 ( .A0(n22486), .A1(sigma12[28]), .B0(n25750), .B1(sigma11[28]), 
        .Y(n24112) );
  NOR2BXL U9455 ( .AN(n4777), .B(n11480), .Y(M3_U3_U1_enc_tree_1__1__28_) );
  AOI22XL U9456 ( .A0(n22486), .A1(sigma12[27]), .B0(n25750), .B1(sigma11[27]), 
        .Y(n25167) );
  AOI22XL U9457 ( .A0(n25763), .A1(n26519), .B0(n25754), .B1(n26455), .Y(
        n25171) );
  AOI22XL U9458 ( .A0(n25763), .A1(n26518), .B0(n25754), .B1(n26448), .Y(
        n24182) );
  NOR2XL U9459 ( .A(M5_a_8_), .B(n15968), .Y(M5_U3_U1_enc_tree_1__1__22_) );
  NOR2XL U9460 ( .A(n5045), .B(n12519), .Y(M3_U3_U1_enc_tree_1__1__18_) );
  INVXL U9461 ( .A(n16869), .Y(n3953) );
  CLKINVX3 U9462 ( .A(n4785), .Y(n16572) );
  AOI22XL U9463 ( .A0(n22486), .A1(sigma12[19]), .B0(n25750), .B1(sigma11[19]), 
        .Y(n24241) );
  NOR2XL U9464 ( .A(n4795), .B(n3022), .Y(M5_U3_U1_enc_tree_1__1__10_) );
  INVXL U9465 ( .A(n12222), .Y(n3736) );
  OR2X1 U9466 ( .A(n25245), .B(n25244), .Y(n23673) );
  INVXL U9467 ( .A(n12595), .Y(n6103) );
  CLKINVX3 U9468 ( .A(n6112), .Y(n18673) );
  NAND2BXL U9469 ( .AN(n16012), .B(n3109), .Y(n4168) );
  NOR2X1 U9470 ( .A(n8112), .B(n8153), .Y(n8156) );
  INVXL U9471 ( .A(n17061), .Y(n5674) );
  NOR2XL U9472 ( .A(M4_a_13_), .B(n18468), .Y(M4_U3_U1_or2_tree_0__1__16_) );
  AOI22XL U9473 ( .A0(n22486), .A1(sigma12[15]), .B0(n25750), .B1(sigma11[15]), 
        .Y(n24207) );
  AOI22XL U9474 ( .A0(n22486), .A1(sigma12[7]), .B0(n25750), .B1(sigma11[7]), 
        .Y(n24146) );
  AOI21XL U9475 ( .A0(M4_a_18_), .A1(n18603), .B0(n3757), .Y(
        M4_U3_U1_enc_tree_0__1__14_) );
  INVXL U9476 ( .A(n16348), .Y(n3623) );
  INVX1 U9477 ( .A(n12758), .Y(n3184) );
  AOI22XL U9478 ( .A0(n22486), .A1(sigma12[13]), .B0(n25750), .B1(sigma11[13]), 
        .Y(n24189) );
  AOI22XL U9479 ( .A0(n25763), .A1(n25917), .B0(n25754), .B1(n26449), .Y(
        n24219) );
  AOI22XL U9480 ( .A0(n22486), .A1(sigma12[0]), .B0(n25750), .B1(sigma11[0]), 
        .Y(n24254) );
  NOR2XL U9481 ( .A(M4_a_9_), .B(n4196), .Y(M4_U3_U1_enc_tree_1__1__22_) );
  AOI22XL U9482 ( .A0(n22486), .A1(sigma12[16]), .B0(n25750), .B1(sigma11[16]), 
        .Y(n24215) );
  CLKINVX3 U9483 ( .A(M3_a_11_), .Y(n12522) );
  NAND2XL U9484 ( .A(n20925), .B(n4875), .Y(n4837) );
  AOI22XL U9485 ( .A0(n25754), .A1(sigma11[21]), .B0(sigma12[21]), .B1(n3059), 
        .Y(n20940) );
  AND2XL U9486 ( .A(n13005), .B(n13004), .Y(n13018) );
  NOR2XL U9487 ( .A(n4888), .B(n18468), .Y(M4_U3_U1_enc_tree_1__1__16_) );
  INVX8 U9488 ( .A(n9087), .Y(n11536) );
  INVXL U9489 ( .A(M3_mult_x_15_b_3_), .Y(n6124) );
  INVX1 U9490 ( .A(n12342), .Y(n3186) );
  INVX4 U9491 ( .A(n9087), .Y(n4566) );
  INVXL U9492 ( .A(n7535), .Y(n5362) );
  INVX1 U9493 ( .A(n18625), .Y(n3187) );
  AOI21XL U9494 ( .A0(n3111), .A1(data[127]), .B0(n4137), .Y(n21168) );
  NAND2XL U9495 ( .A(M3_mult_x_15_b_1_), .B(M3_mult_x_15_b_3_), .Y(n6122) );
  OR2X2 U9496 ( .A(n18168), .B(n18169), .Y(n3407) );
  NOR2X2 U9497 ( .A(n23986), .B(n23985), .Y(n23987) );
  AND2XL U9498 ( .A(n17398), .B(n17397), .Y(n17411) );
  BUFX3 U9499 ( .A(M1_a_10_), .Y(n14118) );
  NOR2X1 U9500 ( .A(n18738), .B(n18737), .Y(n19028) );
  NOR2X1 U9501 ( .A(n14449), .B(n14701), .Y(n14445) );
  XOR2X1 U9502 ( .A(n4888), .B(n18468), .Y(n17491) );
  NOR2X1 U9503 ( .A(n7399), .B(n7839), .Y(n7397) );
  BUFX3 U9504 ( .A(M1_a_16_), .Y(n14266) );
  AND2XL U9505 ( .A(n2993), .B(n14356), .Y(n14358) );
  CLKINVX8 U9506 ( .A(n4195), .Y(n18504) );
  NOR2X1 U9507 ( .A(n17156), .B(n17155), .Y(n17399) );
  OAI22XL U9508 ( .A0(n6319), .A1(n7093), .B0(n7094), .B1(n3603), .Y(n6317) );
  BUFX2 U9509 ( .A(n18141), .Y(n18238) );
  NAND2XL U9510 ( .A(n5363), .B(n5596), .Y(n5359) );
  AND2XL U9511 ( .A(n19027), .B(n19026), .Y(n19040) );
  OR2X2 U9512 ( .A(n7145), .B(n7535), .Y(n5360) );
  INVXL U9513 ( .A(n5067), .Y(n5064) );
  OAI22XL U9514 ( .A0(n6340), .A1(n7094), .B0(n7093), .B1(n3603), .Y(n6310) );
  NAND2X1 U9515 ( .A(n14862), .B(n14903), .Y(n14906) );
  INVXL U9516 ( .A(n4979), .Y(n4431) );
  AOI22XL U9517 ( .A0(n25255), .A1(sigma12[14]), .B0(n3050), .B1(sigma11[14]), 
        .Y(n20734) );
  INVX8 U9518 ( .A(n3257), .Y(n9087) );
  NOR2X1 U9519 ( .A(n11560), .B(n11559), .Y(n13005) );
  XOR2X1 U9520 ( .A(n18169), .B(n3376), .Y(n3230) );
  NAND2BXL U9521 ( .AN(M0_b_2_), .B(n5578), .Y(n5576) );
  NAND2X1 U9522 ( .A(n8098), .B(n8144), .Y(n8112) );
  AND2XL U9523 ( .A(n7534), .B(n5398), .Y(n5397) );
  NAND2X1 U9524 ( .A(n8111), .B(n8150), .Y(n8153) );
  NOR2XL U9525 ( .A(n3529), .B(n7569), .Y(M0_U4_U1_enc_tree_0__1__18_) );
  AOI2BB1XL U9526 ( .A0N(learning_rate[29]), .A1N(n25856), .B0(n24010), .Y(
        n2622) );
  NOR2X1 U9527 ( .A(n11554), .B(n11553), .Y(n13006) );
  INVXL U9528 ( .A(n17832), .Y(n3193) );
  NAND3X1 U9529 ( .A(n11591), .B(n11590), .C(n11589), .Y(n18773) );
  NAND3X1 U9530 ( .A(n11599), .B(n11598), .C(n11597), .Y(n18779) );
  XOR2X1 U9531 ( .A(n4505), .B(n18658), .Y(n17495) );
  XOR2X1 U9532 ( .A(M3_mult_x_15_b_20_), .B(n6014), .Y(n17058) );
  OAI22XL U9533 ( .A0(n25255), .A1(n26139), .B0(n3050), .B1(n26415), .Y(n25209) );
  NOR2X1 U9534 ( .A(n14840), .B(n14883), .Y(n14862) );
  XOR2X1 U9535 ( .A(n6989), .B(n25874), .Y(n6775) );
  NOR2X1 U9536 ( .A(n14861), .B(n14900), .Y(n14903) );
  BUFX3 U9537 ( .A(M1_a_14_), .Y(n14236) );
  NOR2X1 U9538 ( .A(n17162), .B(n17161), .Y(n17398) );
  NOR2X1 U9539 ( .A(n17169), .B(n17168), .Y(n17405) );
  CLKBUFX8 U9540 ( .A(n17501), .Y(n3195) );
  NOR2X1 U9541 ( .A(n19220), .B(n19263), .Y(n19242) );
  BUFX3 U9542 ( .A(M1_a_22_), .Y(n14357) );
  INVXL U9543 ( .A(n13605), .Y(n4254) );
  NOR2X1 U9544 ( .A(n19241), .B(n19282), .Y(n19285) );
  AOI222XL U9545 ( .A0(n23023), .A1(n10749), .B0(n22887), .B1(n3116), .C0(
        n23021), .C1(n22987), .Y(n10761) );
  XOR2X1 U9546 ( .A(n11495), .B(n6014), .Y(n16889) );
  AOI22XL U9547 ( .A0(n25410), .A1(n26536), .B0(n25567), .B1(n26061), .Y(
        n25534) );
  AOI22XL U9548 ( .A0(n25410), .A1(n26534), .B0(n25567), .B1(n26060), .Y(
        n25519) );
  NAND2X1 U9549 ( .A(n19240), .B(n19239), .Y(n19282) );
  AOI22XL U9550 ( .A0(n25815), .A1(y12[24]), .B0(n3050), .B1(y11[24]), .Y(
        n24101) );
  INVX1 U9551 ( .A(M3_a_0_), .Y(n4775) );
  NOR2X1 U9552 ( .A(n18749), .B(n18748), .Y(n19034) );
  AOI22XL U9553 ( .A0(n25786), .A1(n26108), .B0(n25785), .B1(n26454), .Y(
        n25787) );
  AOI22XL U9554 ( .A0(n25025), .A1(y12[28]), .B0(n3050), .B1(y11[28]), .Y(
        n24402) );
  AOI22XL U9555 ( .A0(n25815), .A1(y12[25]), .B0(n3050), .B1(y11[25]), .Y(
        n24356) );
  NAND3X2 U9556 ( .A(n5467), .B(n4397), .C(n4661), .Y(M4_a_9_) );
  NAND2X1 U9557 ( .A(n19231), .B(n19274), .Y(n19241) );
  NOR2X2 U9558 ( .A(n4921), .B(n4920), .Y(n4919) );
  AOI22XL U9559 ( .A0(n25786), .A1(n26107), .B0(n25785), .B1(n26453), .Y(
        n25223) );
  NOR2X1 U9560 ( .A(n7373), .B(n7372), .Y(n7842) );
  NAND2X2 U9561 ( .A(n5988), .B(n5986), .Y(n11485) );
  NAND2X1 U9562 ( .A(n25206), .B(data[102]), .Y(n4532) );
  AOI22XL U9563 ( .A0(n25785), .A1(n26513), .B0(n25786), .B1(n26450), .Y(
        n24265) );
  INVX8 U9564 ( .A(n4796), .Y(n3199) );
  NOR2X1 U9565 ( .A(n7379), .B(n7378), .Y(n7845) );
  NAND3X1 U9566 ( .A(n18758), .B(n18757), .C(n18756), .Y(n19029) );
  AND2XL U9567 ( .A(n4772), .B(data[119]), .Y(n17158) );
  CLKBUFX8 U9568 ( .A(n11484), .Y(M3_mult_x_15_b_21_) );
  NAND2X1 U9569 ( .A(n14851), .B(n14893), .Y(n14861) );
  AOI21X1 U9570 ( .A0(n21291), .A1(n21290), .B0(n21289), .Y(n21392) );
  NAND2X1 U9571 ( .A(n14839), .B(n14881), .Y(n14883) );
  INVXL U9572 ( .A(M4_a_20_), .Y(n4505) );
  NAND3X1 U9573 ( .A(n11579), .B(n11578), .C(n11577), .Y(n18770) );
  INVX1 U9574 ( .A(M0_a_22_), .Y(n6821) );
  NAND3X1 U9575 ( .A(n11583), .B(n11582), .C(n11581), .Y(n18783) );
  NAND2X1 U9576 ( .A(n25206), .B(data[106]), .Y(n4533) );
  INVX1 U9577 ( .A(n25872), .Y(n7827) );
  INVX4 U9578 ( .A(n6324), .Y(n6944) );
  AND2XL U9579 ( .A(n3111), .B(data[120]), .Y(n17161) );
  AND2XL U9580 ( .A(n3111), .B(data[122]), .Y(n17168) );
  NAND3X1 U9581 ( .A(n17172), .B(n17171), .C(n17170), .Y(n17403) );
  NOR2X1 U9582 ( .A(n17175), .B(n17174), .Y(n17402) );
  NAND3X1 U9583 ( .A(n17178), .B(n17177), .C(n17176), .Y(n17400) );
  INVXL U9584 ( .A(n5983), .Y(n5970) );
  NAND2X1 U9585 ( .A(n14860), .B(n14859), .Y(n14900) );
  NOR2X1 U9586 ( .A(n14751), .B(n14812), .Y(n14816) );
  AOI222XL U9587 ( .A0(n22892), .A1(n10775), .B0(n22708), .B1(n10769), .C0(
        n22891), .C1(n23002), .Y(n22732) );
  NAND3X1 U9588 ( .A(n11575), .B(n11574), .C(n11573), .Y(n13007) );
  NAND3X1 U9589 ( .A(n11569), .B(n11568), .C(n11567), .Y(n13010) );
  NOR2X1 U9590 ( .A(n8119), .B(n8048), .Y(n8122) );
  NOR2X1 U9591 ( .A(n11566), .B(n11565), .Y(n13012) );
  NOR2X1 U9592 ( .A(n8017), .B(n8000), .Y(n8020) );
  NAND2X2 U9593 ( .A(n4243), .B(n5891), .Y(M4_a_5_) );
  INVXL U9594 ( .A(n4806), .Y(n5578) );
  NOR2X1 U9595 ( .A(n8141), .B(n8097), .Y(n8144) );
  AND2XL U9596 ( .A(n4772), .B(data[55]), .Y(n11556) );
  NOR2X1 U9597 ( .A(n8128), .B(n8073), .Y(n8131) );
  AND2X2 U9598 ( .A(n9071), .B(n3558), .Y(n3557) );
  NOR2X1 U9599 ( .A(n11572), .B(n11571), .Y(n13009) );
  AND2XL U9600 ( .A(n4772), .B(data[56]), .Y(n11559) );
  NOR2X1 U9601 ( .A(n8110), .B(n8147), .Y(n8111) );
  NAND2X2 U9602 ( .A(n4030), .B(n5872), .Y(M4_a_12_) );
  CLKINVX8 U9603 ( .A(n18169), .Y(n3206) );
  NAND3X1 U9604 ( .A(n4469), .B(n4753), .C(n4754), .Y(n11498) );
  AOI22XL U9605 ( .A0(n25786), .A1(n26369), .B0(n25785), .B1(n25925), .Y(
        n24159) );
  INVX1 U9606 ( .A(M3_mult_x_15_b_2_), .Y(n3208) );
  CLKINVX3 U9607 ( .A(n3117), .Y(n4576) );
  CLKINVX3 U9608 ( .A(n3117), .Y(n4578) );
  CLKINVX3 U9609 ( .A(n3117), .Y(n4577) );
  OR2XL U9610 ( .A(n3115), .B(n23065), .Y(n9155) );
  CLKINVX8 U9611 ( .A(n26488), .Y(n3209) );
  NOR2X1 U9612 ( .A(n8163), .B(n8188), .Y(n8147) );
  INVX8 U9613 ( .A(n16909), .Y(n3211) );
  NAND2X1 U9614 ( .A(n5032), .B(data[74]), .Y(n4398) );
  NOR2XL U9615 ( .A(M0_b_15_), .B(n7621), .Y(M0_U4_U1_enc_tree_1__1__16_) );
  NOR2XL U9616 ( .A(n7569), .B(M0_b_13_), .Y(M0_U4_U1_enc_tree_1__1__18_) );
  NOR2X1 U9617 ( .A(n19271), .B(n19230), .Y(n19274) );
  OR2XL U9618 ( .A(n3115), .B(n21093), .Y(n9144) );
  OR2XL U9619 ( .A(n3115), .B(n23053), .Y(n9151) );
  NOR2X1 U9620 ( .A(n19238), .B(n19277), .Y(n19240) );
  NAND2XL U9621 ( .A(n23023), .B(n22987), .Y(n10767) );
  NAND2XL U9622 ( .A(n25743), .B(y20[21]), .Y(n5558) );
  NAND2XL U9623 ( .A(n25743), .B(y20[19]), .Y(n4814) );
  NOR2BXL U9624 ( .AN(n6476), .B(M0_a_10_), .Y(M0_U3_U1_enc_tree_1__1__20_) );
  NAND2X1 U9625 ( .A(n14750), .B(n14810), .Y(n14812) );
  OAI2BB1X1 U9626 ( .A0N(y10[30]), .A1N(n3224), .B0(n7369), .Y(n7853) );
  NAND2BX2 U9627 ( .AN(n6088), .B(n4014), .Y(M3_a_10_) );
  AOI2BB1X2 U9628 ( .A0N(n25243), .A1N(n23996), .B0(n4465), .Y(n4464) );
  NAND3X1 U9629 ( .A(n7386), .B(n7385), .C(n14416), .Y(n7848) );
  OR2XL U9630 ( .A(n3115), .B(n24006), .Y(n9158) );
  NOR2X1 U9631 ( .A(n14890), .B(n14850), .Y(n14893) );
  NAND3X1 U9632 ( .A(n7381), .B(n7380), .C(n14413), .Y(n7847) );
  NOR2X1 U9633 ( .A(n14856), .B(n14896), .Y(n14860) );
  NOR2X1 U9634 ( .A(n21335), .B(n21385), .Y(n21388) );
  CLKINVX3 U9635 ( .A(M1_b_11_), .Y(n5489) );
  AND2XL U9636 ( .A(n4875), .B(data[58]), .Y(n11565) );
  INVXL U9637 ( .A(M0_a_16_), .Y(n6028) );
  NOR2X1 U9638 ( .A(n19187), .B(n19170), .Y(n19190) );
  OAI2BB1X1 U9639 ( .A0N(y10[29]), .A1N(n3224), .B0(n7390), .Y(n7852) );
  NOR2BX2 U9640 ( .AN(n5347), .B(n4125), .Y(n4124) );
  OAI2BB1XL U9641 ( .A0N(y12[26]), .A1N(n4826), .B0(n9125), .Y(n9128) );
  INVXL U9642 ( .A(n6476), .Y(n7220) );
  OAI21X1 U9643 ( .A0(n6274), .A1(n26217), .B0(n6251), .Y(M0_b_5_) );
  OAI2BB1XL U9644 ( .A0N(y12[28]), .A1N(n4826), .B0(n9132), .Y(n9135) );
  NAND2XL U9645 ( .A(n4139), .B(n4138), .Y(n4137) );
  NAND2XL U9646 ( .A(n23003), .B(n22987), .Y(n22974) );
  OAI21X2 U9647 ( .A0(n7382), .A1(n26004), .B0(n5565), .Y(M0_a_12_) );
  BUFX2 U9648 ( .A(n23154), .Y(n11089) );
  OAI2BB1XL U9649 ( .A0N(y12[23]), .A1N(n4826), .B0(n9114), .Y(n9117) );
  OAI2BB1XL U9650 ( .A0N(y12[24]), .A1N(n4826), .B0(n9118), .Y(n9121) );
  NOR2X1 U9651 ( .A(n14909), .B(n4802), .Y(n14896) );
  NAND2X1 U9652 ( .A(n11546), .B(n11547), .Y(M1_b_22_) );
  INVXL U9653 ( .A(n8423), .Y(n8443) );
  NAND2X2 U9654 ( .A(n6049), .B(n11522), .Y(M1_b_11_) );
  NOR2X1 U9655 ( .A(n14807), .B(n14749), .Y(n14810) );
  INVX1 U9656 ( .A(n8200), .Y(n8135) );
  NOR2X1 U9657 ( .A(n19258), .B(n19218), .Y(n19261) );
  INVX1 U9658 ( .A(n8185), .Y(n8165) );
  INVXL U9659 ( .A(n8478), .Y(n8496) );
  AND2X2 U9660 ( .A(n5294), .B(n11504), .Y(n4478) );
  INVXL U9661 ( .A(n8480), .Y(n8509) );
  CLKINVX3 U9662 ( .A(n4506), .Y(n4225) );
  INVX1 U9663 ( .A(n8181), .Y(n8167) );
  INVXL U9664 ( .A(n8428), .Y(n8474) );
  NOR2X1 U9665 ( .A(n14868), .B(n14826), .Y(n14871) );
  NOR2X2 U9666 ( .A(n5469), .B(n4654), .Y(n17474) );
  INVXL U9667 ( .A(n8425), .Y(n8459) );
  NOR2X1 U9668 ( .A(n19292), .B(n19318), .Y(n19277) );
  NOR2X1 U9669 ( .A(n19248), .B(n19206), .Y(n19251) );
  CLKINVX4 U9670 ( .A(n10770), .Y(n23002) );
  NAND4X1 U9671 ( .A(n7889), .B(n7888), .C(n7887), .D(n7886), .Y(n8193) );
  INVXL U9672 ( .A(n4822), .Y(n6190) );
  NAND4X1 U9673 ( .A(n8090), .B(n8089), .C(n8088), .D(n8087), .Y(n8181) );
  NAND2XL U9674 ( .A(n21166), .B(sigma12[31]), .Y(n4139) );
  OR2X2 U9675 ( .A(n4860), .B(n26369), .Y(n5467) );
  NAND2X1 U9676 ( .A(n17167), .B(n3024), .Y(n20373) );
  NOR2BX2 U9677 ( .AN(n6095), .B(n6094), .Y(n4506) );
  NAND4X1 U9678 ( .A(n8102), .B(n8101), .C(n8100), .D(n8099), .Y(n8185) );
  AOI22X1 U9679 ( .A0(n5480), .A1(sigma10[9]), .B0(in_valid_t), .B1(w2[9]), 
        .Y(n11492) );
  NAND4X1 U9680 ( .A(n8079), .B(n8078), .C(n8077), .D(n8076), .Y(n8200) );
  AOI22X1 U9681 ( .A0(n5480), .A1(sigma11[1]), .B0(w2[33]), .B1(in_valid_t), 
        .Y(n3375) );
  NAND4X1 U9682 ( .A(n8095), .B(n8094), .C(n8093), .D(n8092), .Y(n8208) );
  NAND4X1 U9683 ( .A(n8108), .B(n8107), .C(n8106), .D(n8105), .Y(n8189) );
  NAND4X1 U9684 ( .A(n8064), .B(n8063), .C(n8062), .D(n8061), .Y(n8196) );
  CLKINVX4 U9685 ( .A(n22636), .Y(n23151) );
  NAND2XL U9686 ( .A(n21166), .B(sigma10[23]), .Y(n11555) );
  OR2X2 U9687 ( .A(n19278), .B(n19322), .Y(n19239) );
  INVX1 U9688 ( .A(n14927), .Y(n14913) );
  NAND2X1 U9689 ( .A(n25693), .B(n20748), .Y(n9043) );
  OR2XL U9690 ( .A(n3116), .B(n10749), .Y(n10748) );
  OR2X2 U9691 ( .A(n14923), .B(n14938), .Y(n14859) );
  NAND4X1 U9692 ( .A(n7987), .B(n7986), .C(n7985), .D(n7984), .Y(n8237) );
  NAND4XL U9693 ( .A(n7910), .B(n7909), .C(n7908), .D(n7907), .Y(n8478) );
  NOR2XL U9694 ( .A(n5581), .B(n5580), .Y(n5579) );
  INVXL U9695 ( .A(n19555), .Y(n19583) );
  NAND4X1 U9696 ( .A(n7993), .B(n7992), .C(n7991), .D(n7990), .Y(n8244) );
  AND2X2 U9697 ( .A(n14923), .B(n14938), .Y(n14897) );
  NAND2XL U9698 ( .A(n5480), .B(sigma11[4]), .Y(n5881) );
  NAND2XL U9699 ( .A(n21166), .B(sigma11[28]), .Y(n18753) );
  NAND2XL U9700 ( .A(n5480), .B(sigma11[18]), .Y(n5016) );
  NAND2XL U9701 ( .A(n21166), .B(sigma11[29]), .Y(n18757) );
  NAND2XL U9702 ( .A(n21166), .B(sigma11[30]), .Y(n18736) );
  INVXL U9703 ( .A(n3024), .Y(n4345) );
  NOR2X1 U9704 ( .A(n15440), .B(n14988), .Y(n14807) );
  NAND4XL U9705 ( .A(n7959), .B(n7958), .C(n7957), .D(n7956), .Y(n8254) );
  INVXL U9706 ( .A(n14934), .Y(n14937) );
  INVX1 U9707 ( .A(n19330), .Y(n19265) );
  INVX1 U9708 ( .A(n19326), .Y(n19255) );
  INVXL U9709 ( .A(n19337), .Y(n19340) );
  AOI22XL U9710 ( .A0(n25822), .A1(n25996), .B0(in_valid_w2), .B1(n26417), .Y(
        n25312) );
  INVX1 U9711 ( .A(n19428), .Y(n19932) );
  AOI22XL U9712 ( .A0(n25820), .A1(n26026), .B0(in_valid_w2), .B1(n26418), .Y(
        n25317) );
  INVXL U9713 ( .A(n19318), .Y(n19321) );
  OR2XL U9714 ( .A(n25837), .B(n23789), .Y(n23790) );
  INVXL U9715 ( .A(n4241), .Y(n3861) );
  AOI22XL U9716 ( .A0(n25822), .A1(n26003), .B0(in_valid_w2), .B1(n26432), .Y(
        n25311) );
  INVX1 U9717 ( .A(n19426), .Y(n19927) );
  NOR2XL U9718 ( .A(n4241), .B(n25807), .Y(n3834) );
  INVX1 U9719 ( .A(n19338), .Y(n19299) );
  AOI22XL U9720 ( .A0(n25820), .A1(n26010), .B0(in_valid_w2), .B1(n26420), .Y(
        n25322) );
  AOI22XL U9721 ( .A0(n25822), .A1(n25998), .B0(in_valid_w2), .B1(n26429), .Y(
        n25307) );
  INVX1 U9722 ( .A(n15050), .Y(n15552) );
  AOI22XL U9723 ( .A0(n25822), .A1(n26002), .B0(in_valid_w2), .B1(n26430), .Y(
        n25309) );
  AOI22XL U9724 ( .A0(n25822), .A1(n25999), .B0(in_valid_w2), .B1(n26431), .Y(
        n25310) );
  AOI22XL U9725 ( .A0(n25822), .A1(n25995), .B0(in_valid_w2), .B1(n26433), .Y(
        n25313) );
  AOI22XL U9726 ( .A0(n25820), .A1(n26012), .B0(in_valid_w2), .B1(n26441), .Y(
        n25327) );
  NAND2X1 U9727 ( .A(n3120), .B(y20[31]), .Y(n8218) );
  AOI22XL U9728 ( .A0(n25822), .A1(n26004), .B0(in_valid_w2), .B1(n26435), .Y(
        n25315) );
  AOI22XL U9729 ( .A0(n25820), .A1(n26005), .B0(in_valid_w2), .B1(n26436), .Y(
        n25318) );
  INVXL U9730 ( .A(n14946), .Y(n14949) );
  AOI22XL U9731 ( .A0(n25820), .A1(n26013), .B0(in_valid_w2), .B1(n26419), .Y(
        n25320) );
  AOI22XL U9732 ( .A0(n25820), .A1(n26016), .B0(in_valid_w2), .B1(n26440), .Y(
        n25326) );
  INVX1 U9733 ( .A(n15053), .Y(n15557) );
  INVX1 U9734 ( .A(n15048), .Y(n15547) );
  AOI22XL U9735 ( .A0(n25820), .A1(n26014), .B0(in_valid_w2), .B1(n26437), .Y(
        n25321) );
  NAND2X1 U9736 ( .A(n8104), .B(y20[30]), .Y(n7886) );
  CLKINVX4 U9737 ( .A(n11395), .Y(n3218) );
  INVX1 U9738 ( .A(n14947), .Y(n14875) );
  AOI22XL U9739 ( .A0(n25820), .A1(n26015), .B0(in_valid_w2), .B1(n26438), .Y(
        n25324) );
  AOI22XL U9740 ( .A0(n25820), .A1(n26011), .B0(in_valid_w2), .B1(n26439), .Y(
        n25325) );
  INVX1 U9741 ( .A(n15066), .Y(n15542) );
  BUFX3 U9742 ( .A(n11140), .Y(n11071) );
  INVX1 U9743 ( .A(n14943), .Y(n14919) );
  AOI22XL U9744 ( .A0(n25822), .A1(n26008), .B0(in_valid_w2), .B1(n26434), .Y(
        n25314) );
  INVXL U9745 ( .A(n22867), .Y(n26495) );
  AOI22XL U9746 ( .A0(n25822), .A1(n26000), .B0(in_valid_w2), .B1(n26426), .Y(
        n25304) );
  AOI22XL U9747 ( .A0(n25822), .A1(n26009), .B0(in_valid_w2), .B1(n26424), .Y(
        n25302) );
  AOI22XL U9748 ( .A0(n25822), .A1(n25997), .B0(in_valid_w2), .B1(n26425), .Y(
        n25303) );
  AOI22XL U9749 ( .A0(n25822), .A1(n26001), .B0(in_valid_w2), .B1(n26428), .Y(
        n25306) );
  AOI22XL U9750 ( .A0(n25822), .A1(n26006), .B0(in_valid_w2), .B1(n26427), .Y(
        n25305) );
  AOI22XL U9751 ( .A0(n25822), .A1(n26017), .B0(in_valid_w2), .B1(n26442), .Y(
        n25823) );
  OAI22X1 U9752 ( .A0(n23193), .A1(n25994), .B0(n9107), .B1(n25889), .Y(n11133) );
  OAI211XL U9753 ( .A0(n2972), .A1(iter[0]), .B0(n23985), .C0(n23063), .Y(
        n1750) );
  NOR2XL U9754 ( .A(n23884), .B(n26568), .Y(n4971) );
  NAND2XL U9755 ( .A(n5604), .B(w2[6]), .Y(n5584) );
  NOR2XL U9756 ( .A(n23884), .B(n26550), .Y(n5965) );
  AND2X2 U9757 ( .A(n14427), .B(y10[5]), .Y(n4125) );
  NOR2XL U9758 ( .A(n23884), .B(n26551), .Y(n4810) );
  INVX1 U9759 ( .A(n21414), .Y(n21379) );
  INVX4 U9760 ( .A(n11481), .Y(n11483) );
  NOR2X1 U9761 ( .A(n7382), .B(n26047), .Y(n7383) );
  NAND2XL U9762 ( .A(n25723), .B(temp0[18]), .Y(n4829) );
  NOR2XL U9763 ( .A(n23884), .B(n26549), .Y(n6006) );
  AND2XL U9764 ( .A(temp0[19]), .B(n25723), .Y(n5598) );
  NAND2XL U9765 ( .A(n25723), .B(temp0[4]), .Y(n23472) );
  NAND2XL U9766 ( .A(n4581), .B(n6153), .Y(n6152) );
  NAND2XL U9767 ( .A(n25723), .B(temp0[12]), .Y(n3532) );
  OR2XL U9768 ( .A(n23884), .B(n26562), .Y(n3458) );
  NAND2X1 U9769 ( .A(n14427), .B(y10[9]), .Y(n3285) );
  OAI22XL U9770 ( .A0(n11057), .A1(n25894), .B0(n9107), .B1(n25953), .Y(n11165) );
  NOR2XL U9771 ( .A(n23884), .B(n26521), .Y(n4715) );
  INVX4 U9772 ( .A(n21527), .Y(n3222) );
  NOR2XL U9773 ( .A(n23884), .B(n26531), .Y(n5916) );
  NOR2XL U9774 ( .A(n23884), .B(n26530), .Y(n4241) );
  INVX1 U9775 ( .A(n6274), .Y(n3224) );
  NAND2X1 U9776 ( .A(n6217), .B(y10[31]), .Y(n8221) );
  AOI21X1 U9777 ( .A0(n19349), .A1(n26213), .B0(n8216), .Y(n8217) );
  NAND2X1 U9778 ( .A(n3062), .B(w1[62]), .Y(n7887) );
  AND2XL U9779 ( .A(n21195), .B(n21623), .Y(n21196) );
  AOI22X1 U9780 ( .A0(y11[30]), .A1(n19235), .B0(n19216), .B1(temp2[30]), .Y(
        n19105) );
  AOI22X1 U9781 ( .A0(n3027), .A1(w2[62]), .B0(n3026), .B1(w1[94]), .Y(n19106)
         );
  OR2X2 U9782 ( .A(in_valid_t), .B(n23071), .Y(n23039) );
  NAND2X1 U9783 ( .A(n17167), .B(n23071), .Y(n23133) );
  AOI21X1 U9784 ( .A0(n19349), .A1(n26195), .B0(n19348), .Y(n19350) );
  AOI22X1 U9785 ( .A0(y12[30]), .A1(n19349), .B0(n19216), .B1(temp3[30]), .Y(
        n14858) );
  NAND2XL U9786 ( .A(n2983), .B(temp1[22]), .Y(n6108) );
  NOR2XL U9787 ( .A(n25693), .B(n25963), .Y(n6153) );
  AOI21X1 U9788 ( .A0(n19349), .A1(n26227), .B0(n14964), .Y(n14965) );
  NAND2X1 U9789 ( .A(n3026), .B(w1[63]), .Y(n8219) );
  NAND2XL U9790 ( .A(n10778), .B(n10777), .Y(n11220) );
  NAND2X4 U9791 ( .A(n23997), .B(n26595), .Y(n25059) );
  CLKINVX4 U9792 ( .A(n9108), .Y(n11057) );
  INVX4 U9793 ( .A(n9106), .Y(n9107) );
  NAND2X1 U9794 ( .A(n11178), .B(n11177), .Y(n22716) );
  NAND2X1 U9795 ( .A(n11084), .B(n11083), .Y(n22713) );
  NAND2X1 U9796 ( .A(n21256), .B(w1[30]), .Y(n21327) );
  NOR2X1 U9797 ( .A(in_valid_w2), .B(n21100), .Y(n24015) );
  NAND2XL U9798 ( .A(valid[0]), .B(y10[15]), .Y(n3573) );
  AND2XL U9799 ( .A(n9071), .B(n3556), .Y(n3555) );
  NAND2X1 U9800 ( .A(n23072), .B(n26140), .Y(n7881) );
  AND2X1 U9801 ( .A(n25886), .B(n7885), .Y(n4143) );
  INVX1 U9802 ( .A(n7885), .Y(n23967) );
  AND2X2 U9803 ( .A(n4579), .B(w1[131]), .Y(n4286) );
  MXI2XL U9804 ( .A(data[28]), .B(data[60]), .S0(n3123), .Y(n1642) );
  INVX1 U9805 ( .A(n25151), .Y(n9047) );
  INVXL U9806 ( .A(n25155), .Y(n5240) );
  MXI2XL U9807 ( .A(data[58]), .B(data[90]), .S0(n3123), .Y(n1672) );
  MXI2XL U9808 ( .A(data[24]), .B(data[56]), .S0(n3123), .Y(n1638) );
  MXI2XL U9809 ( .A(data[30]), .B(data[62]), .S0(n3123), .Y(n1644) );
  MXI2XL U9810 ( .A(data[26]), .B(data[58]), .S0(n3123), .Y(n1640) );
  NAND2X1 U9811 ( .A(in_valid_d), .B(w1[139]), .Y(n11522) );
  MXI2XL U9812 ( .A(data[62]), .B(data[94]), .S0(n3123), .Y(n1676) );
  MXI2XL U9813 ( .A(data[87]), .B(data[119]), .S0(n3123), .Y(n1701) );
  NAND2XL U9814 ( .A(in_valid_t), .B(w2[95]), .Y(n4138) );
  NAND2XL U9815 ( .A(in_valid_t), .B(w2[72]), .Y(n5726) );
  INVXL U9816 ( .A(n25898), .Y(n3981) );
  NOR2X2 U9817 ( .A(y11[31]), .B(valid[0]), .Y(n9106) );
  NAND2XL U9818 ( .A(in_valid_t), .B(w2[50]), .Y(n5013) );
  NAND2X1 U9819 ( .A(in_valid_t), .B(w2[49]), .Y(n4669) );
  NOR2XL U9820 ( .A(n15940), .B(n25929), .Y(n3679) );
  INVXL U9821 ( .A(learning_rate[12]), .Y(n23991) );
  NOR2XL U9822 ( .A(n15940), .B(n26000), .Y(n4526) );
  INVXL U9823 ( .A(learning_rate[3]), .Y(n4287) );
  NOR2XL U9824 ( .A(n4581), .B(n26039), .Y(n5580) );
  NAND2X1 U9825 ( .A(in_valid_t), .B(w2[13]), .Y(n4601) );
  NOR2XL U9826 ( .A(n15940), .B(n26002), .Y(n4898) );
  NOR2XL U9827 ( .A(n15940), .B(n25998), .Y(n4963) );
  NOR2XL U9828 ( .A(n15940), .B(n26001), .Y(n4900) );
  NOR2X1 U9829 ( .A(n15940), .B(n26010), .Y(n5418) );
  NAND2XL U9830 ( .A(in_valid_t), .B(w2[91]), .Y(n17170) );
  NAND2XL U9831 ( .A(in_valid_t), .B(learning_rate[26]), .Y(n11589) );
  NOR2XL U9832 ( .A(n15940), .B(n25995), .Y(n6087) );
  NOR2X1 U9833 ( .A(n4583), .B(n6267), .Y(n25154) );
  NOR2X1 U9834 ( .A(n4585), .B(n6255), .Y(n25157) );
  NOR2X1 U9835 ( .A(n4582), .B(n6244), .Y(n25144) );
  NOR2X1 U9836 ( .A(n4582), .B(n6260), .Y(n25142) );
  NOR2X1 U9837 ( .A(n4582), .B(n6233), .Y(n25140) );
  NOR2X1 U9838 ( .A(n4583), .B(n6225), .Y(n25148) );
  INVX1 U9839 ( .A(data_point[7]), .Y(n6246) );
  INVX8 U9840 ( .A(n4586), .Y(n3229) );
  INVX4 U9841 ( .A(in_valid_t), .Y(n17167) );
  NAND2X2 U9842 ( .A(n3230), .B(n18168), .Y(n17937) );
  XOR2X4 U9843 ( .A(n3376), .B(M4_a_1_), .Y(n18168) );
  OAI21X4 U9844 ( .A0(n25796), .A1(n26249), .B0(n3375), .Y(M4_a_1_) );
  OAI21X2 U9845 ( .A0(n25796), .A1(n26267), .B0(n5050), .Y(n3231) );
  NOR2BX4 U9846 ( .AN(n5882), .B(n3232), .Y(n18169) );
  NOR2X4 U9847 ( .A(n18403), .B(n18404), .Y(n18919) );
  NOR2X4 U9848 ( .A(n3321), .B(n3320), .Y(n5232) );
  NOR2X4 U9849 ( .A(n3318), .B(n3319), .Y(n5231) );
  NOR2X4 U9850 ( .A(n3310), .B(n3308), .Y(n5233) );
  NAND3X4 U9851 ( .A(n3236), .B(n4587), .C(n4552), .Y(n20993) );
  NAND4X4 U9852 ( .A(n5233), .B(n5231), .C(n5232), .D(n20642), .Y(n4552) );
  NOR2X4 U9853 ( .A(n3245), .B(n3239), .Y(n10278) );
  OAI21X4 U9854 ( .A0(n3244), .A1(n3243), .B0(n3240), .Y(n3239) );
  AOI21X4 U9855 ( .A0(n3255), .A1(n3249), .B0(n3246), .Y(n3245) );
  NOR2X2 U9856 ( .A(n4141), .B(n3248), .Y(n3247) );
  INVX1 U9857 ( .A(n9832), .Y(n3256) );
  NOR2X4 U9858 ( .A(in_valid_d), .B(n9043), .Y(n3257) );
  OAI21X4 U9859 ( .A0(n10219), .A1(n10217), .B0(n10220), .Y(n10209) );
  NOR2X4 U9860 ( .A(n10131), .B(n10130), .Y(n10219) );
  XNOR2X4 U9861 ( .A(M2_a_8_), .B(M2_a_7_), .Y(n10159) );
  OAI21X4 U9862 ( .A0(n9087), .A1(n25897), .B0(n3258), .Y(M2_a_7_) );
  NOR2X1 U9863 ( .A(n20810), .B(n5306), .Y(n20751) );
  NAND3X4 U9864 ( .A(n23489), .B(n19098), .C(n3260), .Y(n20810) );
  NOR2X2 U9865 ( .A(n19103), .B(n19099), .Y(n3260) );
  NAND2X4 U9866 ( .A(n9055), .B(n3263), .Y(M2_a_3_) );
  NOR2XL U9867 ( .A(n9445), .B(n9383), .Y(n3270) );
  NOR2X1 U9868 ( .A(n9253), .B(n9906), .Y(n3271) );
  XNOR3X2 U9869 ( .A(n10064), .B(n10063), .C(n10062), .Y(n5380) );
  NAND3X1 U9870 ( .A(n5249), .B(n4676), .C(n5248), .Y(n3272) );
  NAND2X4 U9871 ( .A(n4586), .B(n5582), .Y(n6274) );
  NAND2X1 U9872 ( .A(n4121), .B(n17485), .Y(n5306) );
  OAI21X2 U9873 ( .A0(n9739), .A1(n9740), .B0(n9738), .Y(n3281) );
  XNOR2X4 U9874 ( .A(M2_a_10_), .B(n3282), .Y(n10326) );
  NOR2BX4 U9875 ( .AN(n9086), .B(n3283), .Y(n9843) );
  NAND4X4 U9876 ( .A(n4305), .B(n3817), .C(n17483), .D(n17484), .Y(n3308) );
  XOR2X4 U9877 ( .A(n3309), .B(n4665), .Y(n4305) );
  BUFX8 U9878 ( .A(n10403), .Y(n3288) );
  OR2X2 U9879 ( .A(n9209), .B(n10403), .Y(n3289) );
  OR2X2 U9880 ( .A(n9579), .B(n10403), .Y(n3291) );
  OAI22X1 U9881 ( .A0(n4570), .A1(n9218), .B0(n3288), .B1(n9361), .Y(n9339) );
  OAI22X1 U9882 ( .A0(n4570), .A1(n9317), .B0(n3288), .B1(n9297), .Y(n9378) );
  OR2X2 U9883 ( .A(n9617), .B(n3288), .Y(n3294) );
  OR2X2 U9884 ( .A(n10169), .B(n10403), .Y(n3295) );
  OR2X2 U9885 ( .A(n9435), .B(n3288), .Y(n3298) );
  NAND2XL U9886 ( .A(n3299), .B(M2_mult_x_15_n43), .Y(n10454) );
  OAI22X1 U9887 ( .A0(n10367), .A1(n3287), .B0(n3288), .B1(M2_mult_x_15_n43), 
        .Y(n10390) );
  OR2X2 U9888 ( .A(n9651), .B(n3288), .Y(n3300) );
  OR2X2 U9889 ( .A(n9218), .B(n3288), .Y(n3301) );
  NAND2X4 U9890 ( .A(n4365), .B(n4363), .Y(n10635) );
  AOI22X1 U9891 ( .A0(y10[14]), .A1(n14427), .B0(n11536), .B1(n4718), .Y(n5763) );
  NOR2BX4 U9892 ( .AN(n5218), .B(n3307), .Y(n10338) );
  NAND2BX4 U9893 ( .AN(n20269), .B(n17480), .Y(n3310) );
  OAI21X1 U9894 ( .A0(n5237), .A1(n10504), .B0(n10619), .Y(n3311) );
  NAND3X1 U9895 ( .A(n19104), .B(n3050), .C(n20949), .Y(n3314) );
  NAND4BX4 U9896 ( .AN(n10288), .B(n17485), .C(n20711), .D(n20273), .Y(n3319)
         );
  NAND3X2 U9897 ( .A(n5228), .B(n17481), .C(n20808), .Y(n3320) );
  NOR2X1 U9898 ( .A(n3103), .B(n25911), .Y(n5182) );
  NOR2XL U9899 ( .A(n3103), .B(n25916), .Y(n5204) );
  AOI22X2 U9900 ( .A0(n5478), .A1(n23722), .B0(n3128), .B1(n3325), .Y(n25556)
         );
  XOR2X4 U9901 ( .A(n5474), .B(n4701), .Y(n10718) );
  INVX8 U9902 ( .A(n3327), .Y(n14677) );
  NAND2X4 U9903 ( .A(n5276), .B(n5279), .Y(n3327) );
  NAND2X1 U9904 ( .A(n3327), .B(n5501), .Y(n5502) );
  NAND2X1 U9905 ( .A(n3327), .B(n4677), .Y(n4938) );
  NAND2XL U9906 ( .A(n3327), .B(n4561), .Y(n5365) );
  NAND2BXL U9907 ( .AN(n14537), .B(n3327), .Y(n5486) );
  NOR2X1 U9908 ( .A(n3329), .B(n17431), .Y(n3863) );
  NAND2X4 U9909 ( .A(n3331), .B(n3330), .Y(n13898) );
  NAND2X2 U9910 ( .A(n13995), .B(n13994), .Y(n14610) );
  NOR2X4 U9911 ( .A(n13995), .B(n13994), .Y(n14609) );
  NOR2X4 U9912 ( .A(n3332), .B(n3143), .Y(n5211) );
  NOR2X4 U9913 ( .A(n3332), .B(n14724), .Y(n23883) );
  NAND3X4 U9914 ( .A(n4475), .B(n4472), .C(n4474), .Y(n3332) );
  NAND4X4 U9915 ( .A(n17469), .B(n17465), .C(n17423), .D(n17464), .Y(n5699) );
  XNOR3X2 U9916 ( .A(n16019), .B(n16018), .C(n16017), .Y(n6119) );
  NAND2X4 U9917 ( .A(n17147), .B(n15969), .Y(n17148) );
  XOR2X4 U9918 ( .A(n3345), .B(n4590), .Y(n20324) );
  XOR2X4 U9919 ( .A(n3346), .B(n4664), .Y(n3737) );
  XOR2X4 U9920 ( .A(n3348), .B(n4594), .Y(n20970) );
  OAI22X1 U9921 ( .A0(n11783), .A1(n12525), .B0(n12715), .B1(n3350), .Y(n11773) );
  XOR2X1 U9922 ( .A(n5430), .B(n12731), .Y(n3350) );
  NOR2X4 U9923 ( .A(n16856), .B(n16857), .Y(n17220) );
  AND2X4 U9924 ( .A(n3467), .B(n25807), .Y(n23795) );
  NAND2X1 U9925 ( .A(n5312), .B(n3467), .Y(n3462) );
  NOR2X4 U9926 ( .A(n4892), .B(n6106), .Y(n3467) );
  CLKINVX3 U9927 ( .A(n3445), .Y(n3354) );
  NOR2X2 U9928 ( .A(n23519), .B(n3084), .Y(n4201) );
  NOR2XL U9929 ( .A(n23732), .B(n3084), .Y(n23518) );
  CLKINVX8 U9930 ( .A(n5917), .Y(n4220) );
  NAND2X4 U9931 ( .A(n3368), .B(n4023), .Y(n4094) );
  NAND2X2 U9932 ( .A(n4220), .B(n24178), .Y(n4221) );
  NAND2X4 U9933 ( .A(n3355), .B(n18400), .Y(n18918) );
  AOI21X2 U9934 ( .A0(n18791), .A1(n18792), .B0(n3761), .Y(n18833) );
  NAND2BX4 U9935 ( .AN(n18329), .B(n3356), .Y(n18792) );
  NAND2X2 U9936 ( .A(n18330), .B(n18331), .Y(n3356) );
  NAND2X1 U9937 ( .A(n17437), .B(n3357), .Y(n17438) );
  NAND2XL U9938 ( .A(n20346), .B(n3357), .Y(n20347) );
  NAND2XL U9939 ( .A(n20922), .B(n3357), .Y(n20924) );
  OAI21X4 U9940 ( .A0(n3009), .A1(n24262), .B0(n20693), .Y(n3848) );
  INVX8 U9941 ( .A(n21167), .Y(n11479) );
  NAND2X4 U9942 ( .A(n3398), .B(n25693), .Y(n21167) );
  OAI2BB1X4 U9943 ( .A0N(n3365), .A1N(n17210), .B0(n3359), .Y(n3781) );
  AOI2BB1X4 U9944 ( .A0N(n17241), .A1N(n3366), .B0(n3360), .Y(n3359) );
  AOI21X4 U9945 ( .A0(n17216), .A1(n3797), .B0(n3362), .Y(n17241) );
  OAI21X4 U9946 ( .A0(n17229), .A1(n17231), .B0(n17232), .Y(n17216) );
  OAI21X4 U9947 ( .A0(n17204), .A1(n3364), .B0(n3363), .Y(n17210) );
  AOI21X4 U9948 ( .A0(n17205), .A1(n3680), .B0(n5652), .Y(n3363) );
  AOI21X4 U9949 ( .A0(n5656), .A1(n5654), .B0(n5653), .Y(n17204) );
  NAND2X4 U9950 ( .A(n3797), .B(n17249), .Y(n17225) );
  OAI21X2 U9951 ( .A0(n18834), .A1(n18831), .B0(n18835), .Y(n3367) );
  NAND2X1 U9952 ( .A(n18399), .B(n18398), .Y(n18835) );
  NAND2X2 U9953 ( .A(n18397), .B(n18396), .Y(n18831) );
  OAI21X4 U9954 ( .A0(n18731), .A1(n18728), .B0(n18732), .Y(n3761) );
  NOR2X4 U9955 ( .A(n18395), .B(n18394), .Y(n18731) );
  NOR2X4 U9956 ( .A(n18834), .B(n18832), .Y(n4408) );
  NOR2X4 U9957 ( .A(n18397), .B(n18396), .Y(n18832) );
  NOR2X4 U9958 ( .A(n18399), .B(n18398), .Y(n18834) );
  NAND2X4 U9959 ( .A(n5456), .B(n3368), .Y(n3391) );
  NAND3X4 U9960 ( .A(n3839), .B(n3838), .C(n3006), .Y(n3368) );
  NAND2X2 U9961 ( .A(n16855), .B(n16854), .Y(n17253) );
  NOR2X4 U9962 ( .A(n17252), .B(n17220), .Y(n3797) );
  NOR2X2 U9963 ( .A(n16855), .B(n16854), .Y(n17252) );
  OAI22X1 U9964 ( .A0(n17656), .A1(n18242), .B0(n18168), .B1(n3371), .Y(n17697) );
  XNOR2X1 U9965 ( .A(n4206), .B(n3206), .Y(n3413) );
  NAND4X2 U9966 ( .A(n3707), .B(n3787), .C(n3426), .D(n3425), .Y(n3372) );
  NOR2X4 U9967 ( .A(n3699), .B(n3373), .Y(n5335) );
  NOR2X4 U9968 ( .A(n3374), .B(n3862), .Y(n3699) );
  XOR2X4 U9969 ( .A(M5_a_22_), .B(n6014), .Y(n17147) );
  XNOR3X2 U9970 ( .A(n3433), .B(n17545), .C(n17546), .Y(n17652) );
  XNOR3X2 U9971 ( .A(n17534), .B(n5864), .C(n17533), .Y(n3433) );
  OAI22X4 U9972 ( .A0(n17519), .A1(n18242), .B0(n18168), .B1(n3206), .Y(n17534) );
  AOI2BB1X2 U9973 ( .A0N(n3377), .A1N(n3892), .B0(n3891), .Y(n3890) );
  NAND2BX4 U9974 ( .AN(n4415), .B(n4597), .Y(n3725) );
  NOR2X4 U9975 ( .A(n3379), .B(n3378), .Y(n4415) );
  XOR2X4 U9976 ( .A(n3380), .B(n12881), .Y(n23484) );
  AOI2BB1X4 U9977 ( .A0N(n3845), .A1N(n6134), .B0(n12872), .Y(n3380) );
  AOI21X1 U9978 ( .A0(data[33]), .A1(n11479), .B0(n3982), .Y(n3389) );
  INVX2 U9979 ( .A(n3391), .Y(n25128) );
  NAND2X4 U9980 ( .A(n3391), .B(n4698), .Y(n5914) );
  NAND2X2 U9981 ( .A(n3391), .B(n6133), .Y(n6132) );
  NOR2X1 U9982 ( .A(n3391), .B(n20658), .Y(n4174) );
  NOR2XL U9983 ( .A(n3391), .B(n6131), .Y(n6130) );
  NAND2X1 U9984 ( .A(n3391), .B(n6042), .Y(n6041) );
  NAND2XL U9985 ( .A(n3391), .B(n5912), .Y(n3390) );
  CLKINVX4 U9986 ( .A(M4_U3_U1_or2_inv_0__30_), .Y(n18006) );
  NOR2XL U9987 ( .A(n3393), .B(n17432), .Y(n17428) );
  INVX4 U9988 ( .A(n17210), .Y(n17305) );
  NOR2X4 U9989 ( .A(n5639), .B(n3396), .Y(n17038) );
  OAI21X4 U9990 ( .A0(n17213), .A1(n17207), .B0(n17208), .Y(n5652) );
  INVXL U9991 ( .A(n3397), .Y(n18915) );
  NOR2X2 U9992 ( .A(n18907), .B(n3397), .Y(n3830) );
  OAI21X1 U9993 ( .A0(n3397), .A1(n18909), .B0(n18914), .Y(n18409) );
  NOR2X2 U9994 ( .A(n18408), .B(n18407), .Y(n3397) );
  XOR2X4 U9995 ( .A(n3399), .B(n18954), .Y(n23548) );
  XOR2X4 U9996 ( .A(n3400), .B(n4608), .Y(n19019) );
  OAI21X4 U9997 ( .A0(n19014), .A1(n18930), .B0(n18929), .Y(n3400) );
  XOR2X4 U9998 ( .A(n3401), .B(n4593), .Y(n19021) );
  OAI21X4 U9999 ( .A0(n19014), .A1(n18940), .B0(n18939), .Y(n3401) );
  OAI21X1 U10000 ( .A0(n18242), .A1(n3206), .B0(n3407), .Y(n3406) );
  NAND3X1 U10001 ( .A(n5772), .B(n4524), .C(n3411), .Y(n23553) );
  INVXL U10002 ( .A(n20699), .Y(n3411) );
  XOR2X4 U10003 ( .A(n18850), .B(n18849), .Y(n4222) );
  AOI21X4 U10004 ( .A0(n12892), .A1(n3648), .B0(n3647), .Y(n3469) );
  XOR2X4 U10005 ( .A(M4_a_4_), .B(n18169), .Y(n18141) );
  OAI21X1 U10006 ( .A0(n18336), .A1(n18337), .B0(n18335), .Y(n3419) );
  OAI22X2 U10007 ( .A0(n12759), .A1(n11782), .B0(n12760), .B1(n5976), .Y(
        n11891) );
  XOR2X1 U10008 ( .A(n3184), .B(n5430), .Y(n5976) );
  CLKINVX3 U10009 ( .A(n12428), .Y(n3420) );
  NOR2X4 U10010 ( .A(n3423), .B(n17207), .Y(n3680) );
  NOR2X4 U10011 ( .A(n16847), .B(n16846), .Y(n3423) );
  XNOR3X2 U10012 ( .A(n5865), .B(n17609), .C(n17608), .Y(n17648) );
  OAI2BB1X2 U10013 ( .A0N(n4183), .A1N(n17596), .B0(n3428), .Y(n17592) );
  NAND2X2 U10014 ( .A(n18403), .B(n18404), .Y(n18920) );
  INVX8 U10015 ( .A(n3429), .Y(n19014) );
  NAND2BX4 U10016 ( .AN(n18421), .B(n3431), .Y(n3429) );
  INVX1 U10017 ( .A(n3433), .Y(n3432) );
  XOR2X1 U10018 ( .A(n3757), .B(n18467), .Y(n17493) );
  NOR2X4 U10019 ( .A(n3435), .B(n3434), .Y(n18467) );
  NOR2X2 U10020 ( .A(n25796), .B(n26253), .Y(n3434) );
  NOR2X2 U10021 ( .A(n20699), .B(n3014), .Y(n3437) );
  NOR2BX4 U10022 ( .AN(n5464), .B(n23549), .Y(n4508) );
  OAI22X1 U10023 ( .A0(n25813), .A1(n25909), .B0(n24001), .B1(n17167), .Y(
        n3438) );
  NOR2BX1 U10024 ( .AN(n17993), .B(n3439), .Y(n17998) );
  NAND3X2 U10025 ( .A(n20698), .B(n19019), .C(n20701), .Y(n3443) );
  NOR2X4 U10026 ( .A(n3442), .B(n3441), .Y(n3839) );
  NAND3X2 U10027 ( .A(n5637), .B(n23548), .C(n19022), .Y(n3442) );
  NOR2X4 U10028 ( .A(n3444), .B(n3443), .Y(n3838) );
  NAND3X4 U10029 ( .A(n5446), .B(n4185), .C(n4201), .Y(n5033) );
  NOR2X4 U10030 ( .A(n20966), .B(n3446), .Y(n4029) );
  NOR2X4 U10031 ( .A(n12508), .B(n12507), .Y(n12909) );
  NAND2X4 U10032 ( .A(n3137), .B(n4645), .Y(n5985) );
  OAI21X2 U10033 ( .A0(n4597), .A1(n3977), .B0(n3447), .Y(n4645) );
  NAND3X1 U10034 ( .A(n4412), .B(n4415), .C(n4867), .Y(n3447) );
  NAND2X4 U10035 ( .A(n3724), .B(n5932), .Y(n6106) );
  NAND3BX2 U10036 ( .AN(n5400), .B(n12844), .C(n4378), .Y(n3986) );
  NOR2X4 U10037 ( .A(n14614), .B(n14618), .Y(n5210) );
  NOR2X4 U10038 ( .A(n13989), .B(n13990), .Y(n14618) );
  XNOR3X4 U10039 ( .A(n3449), .B(n13825), .C(n13824), .Y(n13990) );
  NOR2X2 U10040 ( .A(n13988), .B(n13987), .Y(n14614) );
  NAND2X2 U10041 ( .A(n3450), .B(n4473), .Y(n4472) );
  NAND4X4 U10042 ( .A(n6073), .B(n14671), .C(n6072), .D(n14670), .Y(n3450) );
  NAND2X4 U10043 ( .A(n4552), .B(n5074), .Y(n5217) );
  NAND2BX4 U10044 ( .AN(n5090), .B(n3454), .Y(n9901) );
  BUFX12 U10045 ( .A(n23892), .Y(n3455) );
  NOR2X4 U10046 ( .A(n4542), .B(n5098), .Y(n23892) );
  AND2X4 U10047 ( .A(n10736), .B(n5097), .Y(n20952) );
  XOR2X4 U10048 ( .A(n3457), .B(n7835), .Y(n10736) );
  OAI21X1 U10049 ( .A0(n3012), .A1(n3605), .B0(n7824), .Y(n3457) );
  AOI21X1 U10050 ( .A0(n3461), .A1(n25796), .B0(n21034), .Y(n2272) );
  INVX1 U10051 ( .A(n3939), .Y(n3466) );
  NAND2XL U10052 ( .A(n3465), .B(n12103), .Y(n3464) );
  OAI21X4 U10053 ( .A0(n3845), .A1(n3719), .B0(n3717), .Y(n12892) );
  NAND3X4 U10054 ( .A(n3726), .B(n3725), .C(n5989), .Y(n4892) );
  XOR2XL U10055 ( .A(n3204), .B(n6162), .Y(n12030) );
  AOI21X4 U10056 ( .A0(n3509), .A1(n3480), .B0(n3479), .Y(n3504) );
  NAND2X4 U10057 ( .A(n5636), .B(n3481), .Y(n3509) );
  NOR2X4 U10058 ( .A(n10736), .B(n3482), .Y(n3604) );
  AOI22X2 U10059 ( .A0(n3483), .A1(n3455), .B0(n20899), .B1(n3139), .Y(n23509)
         );
  NOR2X4 U10060 ( .A(in_valid_d), .B(valid[0]), .Y(n6223) );
  NAND3X4 U10061 ( .A(n3485), .B(n5609), .C(n3484), .Y(n4542) );
  NAND3X2 U10062 ( .A(n5395), .B(n10724), .C(n10727), .Y(n3484) );
  NAND2X2 U10063 ( .A(n3486), .B(n10725), .Y(n3485) );
  CLKINVX4 U10064 ( .A(n5395), .Y(n3486) );
  NAND3X4 U10065 ( .A(n3521), .B(n3487), .C(n3518), .Y(n5395) );
  INVX4 U10066 ( .A(n3524), .Y(n3487) );
  NAND2X1 U10067 ( .A(n3455), .B(n23580), .Y(n3488) );
  NAND2X1 U10068 ( .A(n3455), .B(n20908), .Y(n3490) );
  AOI21X1 U10069 ( .A0(n25738), .A1(n3065), .B0(n4845), .Y(n23902) );
  NAND2X1 U10070 ( .A(n3455), .B(n23893), .Y(n3493) );
  BUFX12 U10071 ( .A(n3605), .Y(n3494) );
  OAI21X2 U10072 ( .A0(n3494), .A1(n7815), .B0(n7822), .Y(n3551) );
  AOI21X4 U10073 ( .A0(n7437), .A1(n3496), .B0(n3495), .Y(n3605) );
  OAI21X4 U10074 ( .A0(n3539), .A1(n7445), .B0(n3606), .Y(n3495) );
  NOR2X4 U10075 ( .A(n3539), .B(n7423), .Y(n3496) );
  OAI21X4 U10076 ( .A0(n7008), .A1(n3583), .B0(n3597), .Y(n7437) );
  NOR2X1 U10077 ( .A(n3500), .B(n25141), .Y(n6236) );
  INVX8 U10078 ( .A(n3499), .Y(n6266) );
  CLKINVX8 U10079 ( .A(n6266), .Y(n6733) );
  NOR2X4 U10080 ( .A(in_valid_d), .B(n3501), .Y(n3499) );
  NOR2X1 U10081 ( .A(n6266), .B(n25894), .Y(n3500) );
  AOI21X4 U10082 ( .A0(n3510), .A1(n3507), .B0(n3503), .Y(n7008) );
  OAI21X4 U10083 ( .A0(n3505), .A1(n3508), .B0(n3504), .Y(n3503) );
  AND2X2 U10084 ( .A(n6723), .B(n6724), .Y(n3506) );
  NOR2X4 U10085 ( .A(n6468), .B(n3508), .Y(n3507) );
  NAND2X4 U10086 ( .A(n3509), .B(n6417), .Y(n3508) );
  NAND2X1 U10087 ( .A(n5555), .B(n5556), .Y(n3514) );
  OAI21X4 U10088 ( .A0(n6274), .A1(n26221), .B0(n6249), .Y(n7569) );
  INVX2 U10089 ( .A(n20760), .Y(n3586) );
  OAI21X2 U10090 ( .A0(n6723), .A1(n6724), .B0(n6728), .Y(n6468) );
  NOR2X4 U10091 ( .A(n3520), .B(n3519), .Y(n3518) );
  NOR2X4 U10092 ( .A(n3523), .B(n3522), .Y(n3521) );
  NAND4BX2 U10093 ( .AN(n3528), .B(n20369), .C(n20832), .D(n20830), .Y(n3524)
         );
  NAND2X1 U10094 ( .A(n10737), .B(n20278), .Y(n3527) );
  OAI21X4 U10095 ( .A0(n26223), .A1(n6274), .B0(n6262), .Y(n7621) );
  XOR2X1 U10096 ( .A(n7073), .B(n7074), .Y(n3533) );
  XOR2X1 U10097 ( .A(n3533), .B(n7075), .Y(n7131) );
  NOR3X4 U10098 ( .A(n20279), .B(n3535), .C(n3534), .Y(n20865) );
  NAND3X1 U10099 ( .A(n3537), .B(n5100), .C(n20283), .Y(n20281) );
  NAND2X4 U10100 ( .A(n7443), .B(n5354), .Y(n3539) );
  NOR2X4 U10101 ( .A(n3546), .B(n3148), .Y(n3545) );
  NAND2BX2 U10102 ( .AN(n20828), .B(n20830), .Y(n3546) );
  AOI21X4 U10103 ( .A0(n3549), .A1(n7321), .B0(n5127), .Y(n7445) );
  NOR2X4 U10104 ( .A(n7308), .B(n7312), .Y(n3549) );
  AOI21XL U10105 ( .A0(n3550), .A1(n25744), .B0(n5557), .Y(n2381) );
  AOI21X1 U10106 ( .A0(n3550), .A1(in_valid_d), .B0(n25729), .Y(n25730) );
  NAND3BX2 U10107 ( .AN(n20755), .B(n20757), .C(n20816), .Y(n20284) );
  NOR2BX4 U10108 ( .AN(n7766), .B(n3553), .Y(n3552) );
  NOR2X4 U10109 ( .A(n3494), .B(n7767), .Y(n3553) );
  NAND2X1 U10110 ( .A(n20762), .B(n20759), .Y(n20755) );
  XOR2X4 U10111 ( .A(n3554), .B(n4609), .Y(n20762) );
  OAI21X2 U10112 ( .A0(n3494), .A1(n7760), .B0(n7759), .Y(n3554) );
  NAND2X1 U10113 ( .A(n7389), .B(y10[19]), .Y(n3559) );
  AOI2BB1X2 U10114 ( .A0N(n6966), .A1N(n7712), .B0(n3565), .Y(n3564) );
  NOR2X1 U10115 ( .A(n6930), .B(n4642), .Y(n3565) );
  INVX2 U10116 ( .A(n7437), .Y(n7446) );
  NAND2BX1 U10117 ( .AN(n7323), .B(n7437), .Y(n3567) );
  XOR2X4 U10118 ( .A(n3571), .B(n7023), .Y(n20951) );
  AOI21X2 U10119 ( .A0(n7364), .A1(n7019), .B0(n7018), .Y(n3571) );
  CLKINVX8 U10120 ( .A(n6266), .Y(n7389) );
  NAND2X4 U10121 ( .A(n3579), .B(n6294), .Y(n7287) );
  NOR2X2 U10122 ( .A(n7268), .B(n7269), .Y(n7438) );
  AOI21X1 U10123 ( .A0(n24743), .A1(n3065), .B0(n23937), .Y(n23938) );
  INVX8 U10124 ( .A(n6223), .Y(n7382) );
  NAND3BX4 U10125 ( .AN(n25147), .B(n3582), .C(n3581), .Y(n4789) );
  NAND2X1 U10126 ( .A(n6223), .B(w2[9]), .Y(n3581) );
  NAND2X1 U10127 ( .A(n6733), .B(y10[9]), .Y(n3582) );
  NAND2X2 U10128 ( .A(n7019), .B(n5099), .Y(n3583) );
  NOR2X4 U10129 ( .A(n7013), .B(n7020), .Y(n5099) );
  NOR2X4 U10130 ( .A(n6910), .B(n6909), .Y(n7020) );
  NOR2X4 U10131 ( .A(n6912), .B(n6911), .Y(n7013) );
  XOR2X1 U10132 ( .A(n6344), .B(n6343), .Y(n6352) );
  INVXL U10133 ( .A(n10741), .Y(n20276) );
  AND2X4 U10134 ( .A(n10741), .B(n10739), .Y(n20855) );
  NOR2X2 U10135 ( .A(n7428), .B(n7446), .Y(n3589) );
  OAI22X1 U10136 ( .A0(n6750), .A1(n6991), .B0(n6990), .B1(n6775), .Y(n6789)
         );
  NAND2X4 U10137 ( .A(n7040), .B(n3590), .Y(n6991) );
  AOI21X4 U10138 ( .A0(n5099), .A1(n7018), .B0(n3592), .Y(n3597) );
  NOR2X4 U10139 ( .A(n6908), .B(n6907), .Y(n7365) );
  INVX1 U10140 ( .A(n6402), .Y(n3594) );
  XNOR2X2 U10141 ( .A(M0_a_4_), .B(M0_a_3_), .Y(n3599) );
  CLKINVX3 U10142 ( .A(n7092), .Y(n26488) );
  NAND2X4 U10143 ( .A(n5620), .B(n6243), .Y(n7092) );
  NAND2X4 U10144 ( .A(n3599), .B(n3598), .Y(n7093) );
  XOR2X1 U10145 ( .A(M0_a_4_), .B(n7092), .Y(n3598) );
  NOR2X4 U10146 ( .A(n4542), .B(n10727), .Y(n10728) );
  OAI21X1 U10147 ( .A0(n3605), .A1(n7487), .B0(n7489), .Y(n7486) );
  AOI21X4 U10148 ( .A0(n7444), .A1(n5354), .B0(n7270), .Y(n3606) );
  OAI22X4 U10149 ( .A0(n3612), .A1(n5655), .B0(n3608), .B1(n3607), .Y(n5653)
         );
  AOI22X1 U10150 ( .A0(n16779), .A1(n16778), .B0(n16781), .B1(n16780), .Y(
        n3607) );
  OAI21X4 U10151 ( .A0(n16778), .A1(n16779), .B0(n3609), .Y(n5655) );
  INVX1 U10152 ( .A(n16781), .Y(n3610) );
  AOI22X2 U10153 ( .A0(n16777), .A1(n3613), .B0(n16775), .B1(n16776), .Y(n3612) );
  AND2X2 U10154 ( .A(n16774), .B(n16773), .Y(n3613) );
  NAND2X4 U10155 ( .A(n16960), .B(n15944), .Y(n16962) );
  OAI22XL U10156 ( .A0(n16962), .A1(n15954), .B0(n16124), .B1(n16960), .Y(
        n16132) );
  OAI21XL U10157 ( .A0(n16103), .A1(n16960), .B0(n3616), .Y(n16441) );
  OAI21XL U10158 ( .A0(n15955), .A1(n16962), .B0(n3617), .Y(n16034) );
  NAND2BXL U10159 ( .AN(n15954), .B(n3637), .Y(n3617) );
  OAI21XL U10160 ( .A0(n16069), .A1(n16962), .B0(n3619), .Y(n16094) );
  OAI21XL U10161 ( .A0(n16069), .A1(n16960), .B0(n3620), .Y(n16796) );
  OAI21XL U10162 ( .A0(n16347), .A1(n16962), .B0(n3621), .Y(n16365) );
  NAND2BXL U10163 ( .AN(n16383), .B(n3637), .Y(n3621) );
  OAI21XL U10164 ( .A0(n16347), .A1(n16960), .B0(n3622), .Y(n16386) );
  XOR2X4 U10165 ( .A(n3199), .B(n5646), .Y(n3637) );
  OAI22X1 U10166 ( .A0(n16883), .A1(n16977), .B0(n3105), .B1(n3199), .Y(n16881) );
  NOR2X1 U10167 ( .A(n15942), .B(n26032), .Y(n3624) );
  NAND2X4 U10168 ( .A(n17427), .B(n3626), .Y(n3852) );
  AOI21X4 U10169 ( .A0(n3085), .A1(n3628), .B0(n3919), .Y(n3626) );
  XOR2X4 U10170 ( .A(n3629), .B(n4702), .Y(n17427) );
  OAI2BB1X4 U10171 ( .A0N(n5339), .A1N(n3781), .B0(n4106), .Y(n3629) );
  OAI2BB1X2 U10172 ( .A0N(n17341), .A1N(n3781), .B0(n17325), .Y(n3932) );
  NAND2XL U10173 ( .A(n3632), .B(n16052), .Y(n3631) );
  NOR2X4 U10174 ( .A(n3893), .B(n4319), .Y(M3_U3_U1_or2_inv_0__18_) );
  CLKINVX3 U10175 ( .A(n3639), .Y(n3638) );
  NAND2X1 U10176 ( .A(n3641), .B(n3640), .Y(n11906) );
  OAI21XL U10177 ( .A0(n11881), .A1(n3114), .B0(n3642), .Y(n3641) );
  OAI22X1 U10178 ( .A0(n12152), .A1(n12265), .B0(n3185), .B1(n4002), .Y(n3642)
         );
  XOR2X1 U10179 ( .A(n11881), .B(n3114), .Y(n3643) );
  XOR3X2 U10180 ( .A(n11716), .B(n11717), .C(n11715), .Y(n11718) );
  NOR2X4 U10181 ( .A(n3646), .B(n4892), .Y(n4950) );
  OAI21X4 U10182 ( .A0(n12891), .A1(n4132), .B0(n3750), .Y(n3647) );
  NOR2X4 U10183 ( .A(n4132), .B(n12890), .Y(n3648) );
  NAND2X4 U10184 ( .A(n12493), .B(n12492), .Y(n3649) );
  NOR2XL U10185 ( .A(n11750), .B(n11751), .Y(n3653) );
  XNOR3X2 U10186 ( .A(n11751), .B(n11750), .C(n3654), .Y(n11840) );
  NOR2X1 U10187 ( .A(n3656), .B(n3655), .Y(n3654) );
  NAND2X2 U10188 ( .A(n4415), .B(n4412), .Y(n3657) );
  NOR2X4 U10189 ( .A(n4414), .B(n4413), .Y(n4412) );
  OAI21X4 U10190 ( .A0(n12907), .A1(n12909), .B0(n12910), .Y(n12902) );
  OAI2BB1X1 U10191 ( .A0N(n11921), .A1N(n3661), .B0(n3659), .Y(n11942) );
  INVXL U10192 ( .A(n3663), .Y(n3660) );
  NAND2XL U10193 ( .A(n3662), .B(n3663), .Y(n3661) );
  XNOR3X2 U10194 ( .A(n3663), .B(n11922), .C(n11921), .Y(n11929) );
  NOR2X1 U10195 ( .A(n11914), .B(n12342), .Y(n3664) );
  INVX1 U10196 ( .A(n11879), .Y(n3665) );
  OAI21X4 U10197 ( .A0(n3415), .A1(n12980), .B0(n3844), .Y(n4367) );
  NAND2X1 U10198 ( .A(n23450), .B(n3668), .Y(n23573) );
  OAI2BB1X1 U10199 ( .A0N(n16514), .A1N(n3671), .B0(n3669), .Y(n16508) );
  NAND2XL U10200 ( .A(n16515), .B(n3670), .Y(n3669) );
  INVXL U10201 ( .A(n3673), .Y(n3670) );
  NAND2BXL U10202 ( .AN(n16515), .B(n3673), .Y(n3671) );
  XOR2X1 U10203 ( .A(n16514), .B(n3672), .Y(n16547) );
  XNOR2X1 U10204 ( .A(n16515), .B(n3673), .Y(n3672) );
  NOR2X1 U10205 ( .A(n3675), .B(n3674), .Y(n3673) );
  NOR2X1 U10206 ( .A(n5835), .B(n16497), .Y(n3674) );
  NOR2XL U10207 ( .A(n16532), .B(n16704), .Y(n3675) );
  NOR2X1 U10208 ( .A(n15940), .B(n25930), .Y(n3677) );
  AOI21X1 U10209 ( .A0(n11479), .A1(data[97]), .B0(n3679), .Y(n3678) );
  OAI22X2 U10210 ( .A0(n16704), .A1(n16116), .B0(n16049), .B1(n5835), .Y(n3686) );
  XOR3X2 U10211 ( .A(n16114), .B(n3686), .C(n16113), .Y(n16813) );
  XOR2X4 U10212 ( .A(n3687), .B(n4604), .Y(n17423) );
  OAI21X2 U10213 ( .A0(n17319), .A1(n3688), .B0(n17324), .Y(n3687) );
  INVXL U10214 ( .A(n16787), .Y(n3690) );
  OAI2BB1X2 U10215 ( .A0N(n3690), .A1N(n3689), .B0(n16785), .Y(n3785) );
  XOR2X1 U10216 ( .A(n4784), .B(n16631), .Y(n15947) );
  XOR2X1 U10217 ( .A(M5_a_2_), .B(n3047), .Y(n15945) );
  NOR2XL U10218 ( .A(M5_mult_x_15_n1), .B(n3047), .Y(
        M5_U3_U1_or2_tree_0__1__28_) );
  NOR2X1 U10219 ( .A(n15942), .B(n26276), .Y(n3691) );
  OAI22X1 U10220 ( .A0(n25796), .A1(n26021), .B0(n25918), .B1(n15940), .Y(
        n3692) );
  XOR2X2 U10221 ( .A(n16090), .B(n3696), .Y(n16789) );
  NOR2X4 U10222 ( .A(n3699), .B(n5658), .Y(n5720) );
  BUFX12 U10223 ( .A(n5720), .Y(n5336) );
  OAI22X1 U10224 ( .A0(n16704), .A1(n16344), .B0(n16343), .B1(n5835), .Y(
        n16357) );
  OAI21X2 U10225 ( .A0(n15997), .A1(n16704), .B0(n3700), .Y(n15991) );
  NAND2BX1 U10226 ( .AN(n15956), .B(n3044), .Y(n3700) );
  NAND2X1 U10227 ( .A(n5847), .B(n2992), .Y(n3701) );
  CLKINVX3 U10228 ( .A(n16704), .Y(n5847) );
  NAND2BX1 U10229 ( .AN(n16380), .B(n3044), .Y(n3702) );
  OAI21X1 U10230 ( .A0(n16434), .A1(n16433), .B0(n16432), .Y(n3703) );
  INVX1 U10231 ( .A(n16433), .Y(n3704) );
  NAND3X1 U10232 ( .A(n3864), .B(n3707), .C(n3863), .Y(n4116) );
  AOI2BB1X4 U10233 ( .A0N(n17204), .A1N(n6144), .B0(n17205), .Y(n3708) );
  XOR2X4 U10234 ( .A(n11485), .B(n5983), .Y(n12342) );
  NAND2BX1 U10235 ( .AN(n12422), .B(n3712), .Y(n3711) );
  XOR2X2 U10236 ( .A(n4013), .B(n12939), .Y(n3713) );
  AOI21X4 U10237 ( .A0(n3715), .A1(n3714), .B0(n3721), .Y(n3845) );
  NOR2X4 U10238 ( .A(n3722), .B(n3716), .Y(n3715) );
  AOI21X4 U10239 ( .A0(n3720), .A1(n12872), .B0(n3718), .Y(n3717) );
  OAI21X4 U10240 ( .A0(n12936), .A1(n12934), .B0(n12937), .Y(n12872) );
  NOR2X4 U10241 ( .A(n12874), .B(n12879), .Y(n3720) );
  OAI21X4 U10242 ( .A0(n3890), .A1(n3722), .B0(n3887), .Y(n3721) );
  OAI21X4 U10243 ( .A0(n12426), .A1(n12425), .B0(n3889), .Y(n3722) );
  NAND3X2 U10244 ( .A(n4412), .B(n24046), .C(n4415), .Y(n3724) );
  OR2X4 U10245 ( .A(n4412), .B(n3723), .Y(n3726) );
  OAI22X1 U10246 ( .A0(n11819), .A1(n12340), .B0(n12338), .B1(n3728), .Y(
        n11818) );
  NAND2BX1 U10247 ( .AN(n11727), .B(n4776), .Y(n3727) );
  XOR2X1 U10248 ( .A(n12446), .B(n12445), .Y(n3729) );
  XOR2X2 U10249 ( .A(n11665), .B(n3733), .Y(n11681) );
  XOR2X1 U10250 ( .A(n11666), .B(n3734), .Y(n3733) );
  OAI21X1 U10251 ( .A0(n11648), .A1(n12352), .B0(n3735), .Y(n3734) );
  OAI22X1 U10252 ( .A0(n11879), .A1(n12342), .B0(n12598), .B1(n3738), .Y(
        n11887) );
  XOR2X1 U10253 ( .A(n3204), .B(n3739), .Y(n3738) );
  INVX1 U10254 ( .A(M3_mult_x_15_b_19_), .Y(n3739) );
  XOR2X1 U10255 ( .A(n11485), .B(n3740), .Y(n11626) );
  NOR2X1 U10256 ( .A(n25796), .B(n26239), .Y(n3741) );
  NAND2X1 U10257 ( .A(n3745), .B(n3743), .Y(n5775) );
  NAND2BX1 U10258 ( .AN(n12446), .B(n11815), .Y(n3744) );
  NOR2X4 U10259 ( .A(n12491), .B(n12490), .Y(n12936) );
  NOR2X4 U10260 ( .A(n12495), .B(n12494), .Y(n12874) );
  NOR2X4 U10261 ( .A(n12493), .B(n12492), .Y(n12879) );
  AOI21X4 U10262 ( .A0(n12926), .A1(n12504), .B0(n3746), .Y(n12891) );
  OAI21X2 U10263 ( .A0(n12886), .A1(n12931), .B0(n12887), .Y(n3746) );
  NOR2X4 U10264 ( .A(n12501), .B(n12500), .Y(n12930) );
  NOR2X4 U10265 ( .A(n12503), .B(n12502), .Y(n12886) );
  OAI21X4 U10266 ( .A0(n12897), .A1(n12895), .B0(n12898), .Y(n12926) );
  NAND2X2 U10267 ( .A(n12499), .B(n12498), .Y(n12898) );
  NOR2X4 U10268 ( .A(n12499), .B(n12498), .Y(n12897) );
  OAI21X1 U10269 ( .A0(n11785), .A1(n4863), .B0(n11784), .Y(n4862) );
  INVX4 U10270 ( .A(n3747), .Y(n5989) );
  NOR2X2 U10271 ( .A(n3748), .B(n3747), .Y(n23485) );
  NAND3X4 U10272 ( .A(n3842), .B(n3843), .C(n3984), .Y(n3747) );
  INVX4 U10273 ( .A(n3749), .Y(n3894) );
  NOR2X1 U10274 ( .A(n3749), .B(n20307), .Y(n20308) );
  NOR2X1 U10275 ( .A(n3749), .B(n23651), .Y(n20311) );
  NOR2X1 U10276 ( .A(n21044), .B(n3749), .Y(n21045) );
  NOR2X1 U10277 ( .A(n4042), .B(n3749), .Y(n4902) );
  NAND2X4 U10278 ( .A(n3910), .B(n3909), .Y(n3749) );
  AOI21X4 U10279 ( .A0(n12902), .A1(n4948), .B0(n4947), .Y(n3750) );
  NAND2X1 U10280 ( .A(n25128), .B(n24110), .Y(n6031) );
  XNOR2X1 U10281 ( .A(n17774), .B(n17772), .Y(n3751) );
  OAI22XL U10282 ( .A0(n12717), .A1(n3754), .B0(n12005), .B1(n12718), .Y(
        n12037) );
  INVX1 U10283 ( .A(n12716), .Y(n3755) );
  NOR4X2 U10284 ( .A(n21037), .B(n3911), .C(n3144), .D(n4001), .Y(n3759) );
  NAND3X2 U10285 ( .A(n3145), .B(n13029), .C(n13028), .Y(n3911) );
  NOR2X1 U10286 ( .A(n17457), .B(n13038), .Y(n3760) );
  INVXL U10287 ( .A(n3766), .Y(n3765) );
  XNOR3X2 U10288 ( .A(n3766), .B(n17720), .C(n17719), .Y(n18363) );
  NOR2X1 U10289 ( .A(n3768), .B(n3767), .Y(n3766) );
  NOR2X1 U10290 ( .A(n17718), .B(n17937), .Y(n3767) );
  NOR2XL U10291 ( .A(n17656), .B(n18168), .Y(n3768) );
  CLKINVX4 U10292 ( .A(n6132), .Y(n25127) );
  NAND2X1 U10293 ( .A(n3773), .B(n6132), .Y(n3772) );
  NAND2X1 U10294 ( .A(n25128), .B(n20787), .Y(n3773) );
  XOR2X1 U10295 ( .A(n16829), .B(n16828), .Y(n3775) );
  NAND2X1 U10296 ( .A(n3777), .B(n3776), .Y(n16833) );
  NAND2XL U10297 ( .A(n16819), .B(n16820), .Y(n3776) );
  OR2X2 U10298 ( .A(n16819), .B(n16820), .Y(n3778) );
  XNOR3X2 U10299 ( .A(n3779), .B(n16818), .C(n16819), .Y(n16841) );
  OAI21X4 U10300 ( .A0(n17260), .A1(n17258), .B0(n17261), .Y(n17205) );
  NOR2X4 U10301 ( .A(n16845), .B(n16844), .Y(n17260) );
  OAI22X1 U10302 ( .A0(n3102), .A1(n16331), .B0(n16332), .B1(n3780), .Y(n16445) );
  XNOR2X1 U10303 ( .A(n12701), .B(n16289), .Y(n3780) );
  NOR2X1 U10304 ( .A(n17371), .B(n17309), .Y(n17353) );
  NAND2X2 U10305 ( .A(n17124), .B(n17311), .Y(n17371) );
  NOR2X4 U10306 ( .A(n16849), .B(n16848), .Y(n17207) );
  NAND2BX1 U10307 ( .AN(n17330), .B(n3781), .Y(n4131) );
  NAND2XL U10308 ( .A(n3781), .B(n3149), .Y(n3808) );
  NAND2BXL U10309 ( .AN(n17357), .B(n3781), .Y(n3786) );
  AOI21X1 U10310 ( .A0(n17377), .A1(n3781), .B0(n17381), .Y(n5650) );
  XOR2X1 U10311 ( .A(n3781), .B(n4646), .Y(n5834) );
  AND2X2 U10312 ( .A(n3781), .B(n17347), .Y(n3793) );
  XNOR2XL U10313 ( .A(M3_mult_x_15_b_13_), .B(n3203), .Y(n15973) );
  OAI22X1 U10314 ( .A0(n16317), .A1(n15972), .B0(n16064), .B1(n17092), .Y(
        n16014) );
  NAND2X4 U10315 ( .A(n17099), .B(n15951), .Y(n17092) );
  NAND2X1 U10316 ( .A(n3785), .B(n3784), .Y(n16084) );
  NAND2XL U10317 ( .A(n16787), .B(n16786), .Y(n3784) );
  NOR2X1 U10318 ( .A(n16766), .B(n3788), .Y(n16567) );
  INVXL U10319 ( .A(n16638), .Y(n3790) );
  OAI21XL U10320 ( .A0(n16684), .A1(n16638), .B0(n3791), .Y(n16542) );
  XNOR2X2 U10321 ( .A(M5_a_10_), .B(n15968), .Y(n15949) );
  XNOR2X1 U10322 ( .A(n16873), .B(M5_a_10_), .Y(n3796) );
  NAND2X1 U10323 ( .A(n16169), .B(n16170), .Y(n3798) );
  XOR3X2 U10324 ( .A(n16170), .B(n16169), .C(n3800), .Y(n16188) );
  OAI21X2 U10325 ( .A0(n4129), .A1(n16151), .B0(n16150), .Y(n3801) );
  OAI22XL U10326 ( .A0(n3102), .A1(n15959), .B0(n16332), .B1(n3802), .Y(n16031) );
  OAI22X1 U10327 ( .A0(n3102), .A1(n3802), .B0(n16332), .B1(n4126), .Y(n16134)
         );
  XOR2XL U10328 ( .A(n16289), .B(n5718), .Y(n3802) );
  NAND2X1 U10329 ( .A(n17375), .B(n3808), .Y(n3807) );
  OAI22XL U10330 ( .A0(n3810), .A1(n16688), .B0(n16126), .B1(n16942), .Y(
        n16176) );
  OAI22XL U10331 ( .A0(n4177), .A1(n16943), .B0(n3810), .B1(n16942), .Y(n16207) );
  XOR2XL U10332 ( .A(n15968), .B(n5718), .Y(n3810) );
  OAI21X1 U10333 ( .A0(n16187), .A1(n3814), .B0(n16186), .Y(n3811) );
  INVX1 U10334 ( .A(n16187), .Y(n3812) );
  NOR2X2 U10335 ( .A(n5320), .B(n23533), .Y(n5319) );
  AOI21XL U10336 ( .A0(n24633), .A1(n24525), .B0(n3819), .Y(n2466) );
  OAI21XL U10337 ( .A0(n17632), .A1(n3823), .B0(n17631), .Y(n3822) );
  INVXL U10338 ( .A(n3824), .Y(n3823) );
  XNOR3X2 U10339 ( .A(n3824), .B(n17631), .C(n17632), .Y(n17611) );
  NOR2X1 U10340 ( .A(n3826), .B(n3825), .Y(n3824) );
  NOR2X1 U10341 ( .A(n17619), .B(n18625), .Y(n3825) );
  NOR2X1 U10342 ( .A(n17506), .B(n18624), .Y(n3826) );
  NOR2BXL U10343 ( .AN(n10338), .B(M2_a_12_), .Y(M2_U3_U1_enc_tree_1__1__18_)
         );
  NOR2XL U10344 ( .A(M2_mult_x_15_n43), .B(n3827), .Y(
        M2_U3_U1_or2_tree_0__1__16_) );
  XOR2X1 U10345 ( .A(M2_a_14_), .B(n10338), .Y(n4559) );
  XOR2X4 U10346 ( .A(n5761), .B(n3827), .Y(n10403) );
  CLKINVX3 U10347 ( .A(n10338), .Y(n3827) );
  OAI21X2 U10348 ( .A0(n10213), .A1(n10244), .B0(n10214), .Y(n5236) );
  NAND2X1 U10349 ( .A(n10134), .B(n3828), .Y(n10214) );
  XOR3X4 U10350 ( .A(n4304), .B(n9268), .C(n9369), .Y(n10133) );
  XOR2X2 U10351 ( .A(n4176), .B(n9368), .Y(n4304) );
  NOR2X4 U10352 ( .A(n10134), .B(n3828), .Y(n10213) );
  NAND2X1 U10353 ( .A(n3830), .B(n18903), .Y(n4170) );
  AOI21X2 U10354 ( .A0(n3830), .A1(n18904), .B0(n18409), .Y(n18866) );
  OAI22X1 U10355 ( .A0(n9264), .A1(n10368), .B0(n10369), .B1(n3831), .Y(n9213)
         );
  XNOR2X1 U10356 ( .A(n10339), .B(n10337), .Y(n3831) );
  OAI22X1 U10357 ( .A0(n25483), .A1(n4583), .B0(n3834), .B1(n3832), .Y(n2593)
         );
  NAND3X1 U10358 ( .A(n4223), .B(n4221), .C(n3861), .Y(n3833) );
  NAND2X2 U10359 ( .A(n24179), .B(n4215), .Y(n4223) );
  OAI21XL U10360 ( .A0(n17643), .A1(n17644), .B0(n17642), .Y(n3836) );
  NAND4X4 U10361 ( .A(n3839), .B(n3838), .C(n3006), .D(n20655), .Y(n5438) );
  XOR2X4 U10362 ( .A(n4777), .B(n2980), .Y(n12284) );
  NAND2X1 U10363 ( .A(n21166), .B(n3981), .Y(n3840) );
  AND2X4 U10364 ( .A(n4525), .B(n4528), .Y(n4777) );
  INVX12 U10365 ( .A(M5_a_0_), .Y(n16475) );
  XNOR3X2 U10366 ( .A(n4075), .B(n3175), .C(n12631), .Y(n12652) );
  OAI22X1 U10367 ( .A0(n12592), .A1(n3841), .B0(n12717), .B1(n12593), .Y(n5414) );
  NAND2X1 U10368 ( .A(n4003), .B(n4700), .Y(n3842) );
  OAI21X2 U10369 ( .A0(n16416), .A1(n16417), .B0(n16415), .Y(n5853) );
  NAND2X4 U10370 ( .A(n12763), .B(n12764), .Y(n3844) );
  AOI2BB1X1 U10371 ( .A0N(n3845), .A1N(n12933), .B0(n12935), .Y(n4013) );
  AOI21X1 U10372 ( .A0(n12865), .A1(n12984), .B0(n12989), .Y(n12797) );
  XOR3X2 U10373 ( .A(n4129), .B(n16151), .C(n16150), .Y(n16154) );
  XOR2X2 U10374 ( .A(n3847), .B(n16147), .Y(n4129) );
  NOR2XL U10375 ( .A(n17427), .B(n3850), .Y(n24260) );
  XNOR2X1 U10376 ( .A(n17966), .B(n3857), .Y(n3856) );
  NOR2X1 U10377 ( .A(n18625), .B(n3207), .Y(n3857) );
  NAND2X4 U10378 ( .A(n15945), .B(n5835), .Y(n16704) );
  NAND2X2 U10379 ( .A(n16860), .B(n16861), .Y(n17300) );
  NOR2X4 U10380 ( .A(n16860), .B(n16861), .Y(n17299) );
  XOR2X1 U10381 ( .A(n3107), .B(n12233), .Y(n6105) );
  XOR2X1 U10382 ( .A(n3199), .B(n3107), .Y(n5037) );
  NAND2BX4 U10383 ( .AN(n3865), .B(n4094), .Y(n19043) );
  NAND2X2 U10384 ( .A(n4244), .B(n5438), .Y(n3865) );
  NAND2XL U10385 ( .A(n3870), .B(n3869), .Y(n3868) );
  XNOR3X2 U10386 ( .A(n17706), .B(n3870), .C(n17705), .Y(n18361) );
  CLKINVX3 U10387 ( .A(M4_a_1_), .Y(M4_U3_U1_or2_inv_0__30_) );
  OAI21X4 U10388 ( .A0(n23436), .A1(n23486), .B0(n23437), .Y(n3938) );
  NAND2X2 U10389 ( .A(n3871), .B(n4986), .Y(n23437) );
  NOR2X4 U10390 ( .A(n5989), .B(n3983), .Y(n3871) );
  OAI21XL U10391 ( .A0(n12100), .A1(n12618), .B0(n3872), .Y(n12096) );
  INVX1 U10392 ( .A(n12271), .Y(n3876) );
  NOR2X1 U10393 ( .A(n23748), .B(n3878), .Y(n3877) );
  NAND2X1 U10394 ( .A(n3895), .B(n13037), .Y(n3878) );
  CLKINVX3 U10395 ( .A(n20668), .Y(n5978) );
  NAND2XL U10396 ( .A(n3882), .B(n25807), .Y(n4952) );
  NOR2X4 U10397 ( .A(n12906), .B(n12909), .Y(n12901) );
  AOI2BB2X2 U10398 ( .B0(n4991), .B1(n4968), .A0N(n12616), .A1N(n3883), .Y(
        n4990) );
  OAI2BB1X2 U10399 ( .A0N(n5973), .A1N(n11873), .B0(n5972), .Y(n4974) );
  INVX4 U10400 ( .A(n12892), .Y(n12929) );
  AOI21X1 U10401 ( .A0(n12892), .A1(n3153), .B0(n3886), .Y(n3885) );
  AND2X2 U10402 ( .A(n12425), .B(n12426), .Y(n3888) );
  AND2X2 U10403 ( .A(n12423), .B(n12424), .Y(n3891) );
  NAND2X1 U10404 ( .A(n12421), .B(n12422), .Y(n3892) );
  NAND2X4 U10405 ( .A(n5942), .B(n12616), .Y(n12618) );
  AOI21X1 U10406 ( .A0(n3894), .A1(n3895), .B0(n13038), .Y(n4052) );
  XNOR3X2 U10407 ( .A(n11752), .B(n3902), .C(n3899), .Y(n11861) );
  NOR2X1 U10408 ( .A(n11790), .B(n11791), .Y(n3901) );
  NOR2XL U10409 ( .A(M3_mult_x_15_a_15_), .B(n12519), .Y(
        M3_U3_U1_or2_tree_0__1__16_) );
  XOR2XL U10410 ( .A(M3_mult_x_15_b_19_), .B(n3903), .Y(n11980) );
  XOR2XL U10411 ( .A(M5_b_18_), .B(n3903), .Y(n11951) );
  XOR2X1 U10412 ( .A(n3021), .B(n3903), .Y(n11878) );
  XOR2X1 U10413 ( .A(n12803), .B(n3903), .Y(n12632) );
  XNOR2XL U10414 ( .A(n6112), .B(n3903), .Y(n12634) );
  XOR2X1 U10415 ( .A(n3201), .B(n3903), .Y(n11915) );
  XOR2X1 U10416 ( .A(n3106), .B(n12519), .Y(n6040) );
  INVX1 U10417 ( .A(n21037), .Y(n23450) );
  NAND2X4 U10418 ( .A(n4029), .B(n20967), .Y(n21037) );
  NOR2X4 U10419 ( .A(n21022), .B(n4028), .Y(n20967) );
  NOR2X4 U10420 ( .A(n12905), .B(n12922), .Y(n4948) );
  NOR2X4 U10421 ( .A(n12512), .B(n12511), .Y(n12922) );
  MXI2X1 U10422 ( .A(mul5_out[15]), .B(n5948), .S0(n5032), .Y(n2326) );
  NAND2X1 U10423 ( .A(n4866), .B(n5949), .Y(mul5_out[15]) );
  XOR2X2 U10424 ( .A(n11974), .B(n3923), .Y(n11972) );
  XOR2X1 U10425 ( .A(n11975), .B(n3924), .Y(n3923) );
  INVX1 U10426 ( .A(n11977), .Y(n3925) );
  XOR3X2 U10427 ( .A(n11833), .B(n3929), .C(n11832), .Y(n12443) );
  OAI21X2 U10428 ( .A0(n12357), .A1(n11794), .B0(n4135), .Y(n3929) );
  NAND2X1 U10429 ( .A(n4382), .B(n3131), .Y(n5952) );
  OAI22X1 U10430 ( .A0(n12759), .A1(n3930), .B0(n11984), .B1(n12760), .Y(n5373) );
  OAI22X1 U10431 ( .A0(n11917), .A1(n12759), .B0(n12760), .B1(n3930), .Y(
        n11955) );
  XOR2X1 U10432 ( .A(n16884), .B(n3184), .Y(n3930) );
  NAND4X1 U10433 ( .A(n5834), .B(n20739), .C(n17445), .D(n17413), .Y(n3934) );
  OAI22X1 U10434 ( .A0(n16638), .A1(n3935), .B0(n16335), .B1(n16475), .Y(
        n16339) );
  NAND2XL U10435 ( .A(n3937), .B(n3109), .Y(n3936) );
  XOR2X1 U10436 ( .A(M5_mult_x_15_n1), .B(n3201), .Y(n3937) );
  XNOR2X1 U10437 ( .A(n4777), .B(n11480), .Y(n11624) );
  OAI22XL U10438 ( .A0(n16238), .A1(n16688), .B0(n4177), .B1(n16942), .Y(
        n16248) );
  NAND2X4 U10439 ( .A(n15967), .B(n16943), .Y(n16942) );
  INVXL U10440 ( .A(n3938), .Y(n5403) );
  INVXL U10441 ( .A(n12104), .Y(n3940) );
  OAI22X1 U10442 ( .A0(n3183), .A1(n12010), .B0(n12357), .B1(n3941), .Y(n12068) );
  XNOR2X1 U10443 ( .A(n12282), .B(n12701), .Y(n3941) );
  AOI21X1 U10444 ( .A0(n3943), .A1(n16770), .B0(n16769), .Y(n16771) );
  NAND2BX1 U10445 ( .AN(n16768), .B(n3942), .Y(n16770) );
  NOR3X2 U10446 ( .A(n17200), .B(n23634), .C(n25136), .Y(n17265) );
  AOI21X1 U10447 ( .A0(n17327), .A1(n17331), .B0(n17114), .Y(n17320) );
  OAI2BB1X2 U10448 ( .A0N(n5336), .A1N(n20742), .B0(n3950), .Y(mul5_out[7]) );
  NAND3X4 U10449 ( .A(n4102), .B(n4103), .C(n17123), .Y(n5667) );
  NAND2X1 U10450 ( .A(n17108), .B(n17109), .Y(n17317) );
  INVX1 U10451 ( .A(n20929), .Y(n3957) );
  NOR2X1 U10452 ( .A(n3958), .B(n20929), .Y(n4653) );
  NAND3BX2 U10453 ( .AN(n17441), .B(n17445), .C(n17443), .Y(n5714) );
  XOR2X4 U10454 ( .A(n3959), .B(n17308), .Y(n17443) );
  NAND2X1 U10455 ( .A(n20739), .B(n17455), .Y(n17441) );
  XOR2X4 U10456 ( .A(n3960), .B(n17302), .Y(n20739) );
  OAI22X1 U10457 ( .A0(n16962), .A1(n16183), .B0(n16960), .B1(n3961), .Y(
        n16218) );
  OAI22X1 U10458 ( .A0(n16962), .A1(n3961), .B0(n16960), .B1(n16239), .Y(
        n16237) );
  XNOR2X1 U10459 ( .A(n12701), .B(n3211), .Y(n3961) );
  NAND2X1 U10460 ( .A(n17236), .B(n3161), .Y(n17242) );
  NOR2X4 U10461 ( .A(n17299), .B(n17227), .Y(n17236) );
  NAND3X1 U10462 ( .A(n23632), .B(n3963), .C(n3962), .Y(n2544) );
  NAND2BX1 U10463 ( .AN(n24626), .B(n3229), .Y(n3962) );
  AOI22XL U10464 ( .A0(n24169), .A1(n23795), .B0(n2984), .B1(temp1[10]), .Y(
        n3963) );
  NAND2X4 U10465 ( .A(n12521), .B(n3112), .Y(n12535) );
  XOR2X4 U10466 ( .A(M3_mult_x_15_n61), .B(n3112), .Y(n12521) );
  OAI22X1 U10467 ( .A0(n12535), .A1(n3021), .B0(n12995), .B1(
        M3_mult_x_15_b_17_), .Y(n3969) );
  NOR2X1 U10468 ( .A(n12782), .B(n12781), .Y(n12866) );
  NAND2XL U10469 ( .A(n3976), .B(n23794), .Y(n23713) );
  NAND2XL U10470 ( .A(n3976), .B(n25329), .Y(n3975) );
  XOR3X2 U10471 ( .A(n12677), .B(n12675), .C(n12676), .Y(n12681) );
  INVX8 U10472 ( .A(n21166), .Y(n15942) );
  OAI21X4 U10473 ( .A0(n13036), .A1(n13035), .B0(n23484), .Y(n3983) );
  NAND2X1 U10474 ( .A(n5400), .B(n3988), .Y(n3987) );
  NOR2X1 U10475 ( .A(n4378), .B(n12844), .Y(n3989) );
  NAND3X2 U10476 ( .A(n20670), .B(n13027), .C(n20671), .Y(n20668) );
  XNOR2X4 U10477 ( .A(n3990), .B(n4627), .Y(n13027) );
  OAI21X4 U10478 ( .A0(n3415), .A1(n12985), .B0(n4080), .Y(n3990) );
  OAI21X1 U10479 ( .A0(n3994), .A1(n3993), .B0(n3991), .Y(n12179) );
  OAI21XL U10480 ( .A0(n12185), .A1(n3992), .B0(n12184), .Y(n3991) );
  INVXL U10481 ( .A(n3994), .Y(n3992) );
  XNOR3X2 U10482 ( .A(n3994), .B(n12185), .C(n12184), .Y(n12211) );
  NOR2X1 U10483 ( .A(n3996), .B(n3995), .Y(n3994) );
  NOR2XL U10484 ( .A(n12173), .B(n12025), .Y(n3995) );
  NOR2X1 U10485 ( .A(n3183), .B(n12150), .Y(n3996) );
  NAND2X1 U10486 ( .A(n4504), .B(n3186), .Y(n6009) );
  NAND2X1 U10487 ( .A(n13024), .B(n21043), .Y(n4001) );
  NOR2XL U10488 ( .A(n12265), .B(n11485), .Y(M3_U3_U1_or2_tree_0__1__24_) );
  XNOR2X4 U10489 ( .A(n4434), .B(n4002), .Y(n12222) );
  AND2X4 U10490 ( .A(n4962), .B(n4964), .Y(n4002) );
  OAI21XL U10491 ( .A0(n3185), .A1(n4008), .B0(n4006), .Y(n12168) );
  OR2XL U10492 ( .A(n12151), .B(n12152), .Y(n4006) );
  OR2XL U10493 ( .A(n12117), .B(n3185), .Y(n4007) );
  XNOR2X1 U10494 ( .A(n12265), .B(n16884), .Y(n4008) );
  NOR2X1 U10495 ( .A(n25328), .B(n4009), .Y(n24240) );
  NAND3X1 U10496 ( .A(n3894), .B(n5978), .C(n3895), .Y(n4010) );
  INVX8 U10497 ( .A(n11479), .Y(n25813) );
  AOI21X1 U10498 ( .A0(data[42]), .A1(n11479), .B0(n6087), .Y(n4014) );
  XNOR2XL U10499 ( .A(n12594), .B(M3_mult_x_15_b_13_), .Y(n11674) );
  OAI21X4 U10500 ( .A0(n25813), .A1(n26235), .B0(n11490), .Y(
        M3_mult_x_15_b_13_) );
  OAI21XL U10501 ( .A0(n12215), .A1(n4019), .B0(n12214), .Y(n4015) );
  OAI22X1 U10502 ( .A0(n12120), .A1(n12338), .B0(n12340), .B1(n4022), .Y(
        n12148) );
  OAI22XL U10503 ( .A0(n12170), .A1(n12340), .B0(n12338), .B1(n4022), .Y(n5509) );
  XOR2X1 U10504 ( .A(n12560), .B(n4239), .Y(n4022) );
  OAI22X1 U10505 ( .A0(n18083), .A1(n17671), .B0(n18429), .B1(n4027), .Y(
        n17676) );
  OAI22X2 U10506 ( .A0(n18083), .A1(n4027), .B0(n18429), .B1(n17539), .Y(n5923) );
  XOR2X2 U10507 ( .A(n12561), .B(n18428), .Y(n4027) );
  NOR2BX1 U10508 ( .AN(n24192), .B(n25328), .Y(n24195) );
  OAI22X1 U10509 ( .A0(n12597), .A1(n11674), .B0(n11650), .B1(n12523), .Y(
        n4751) );
  XNOR2X1 U10510 ( .A(n12701), .B(n12594), .Y(n11650) );
  NAND2X2 U10511 ( .A(n21019), .B(n21017), .Y(n4028) );
  NOR2X1 U10512 ( .A(n3093), .B(n3097), .Y(n4668) );
  AOI22X1 U10513 ( .A0(n5770), .A1(data[76]), .B0(w2[44]), .B1(in_valid_t), 
        .Y(n4030) );
  OAI21XL U10514 ( .A0(n17763), .A1(n17764), .B0(n17762), .Y(n17766) );
  AOI2BB1X2 U10515 ( .A0N(n21029), .A1N(n4772), .B0(n21028), .Y(n2270) );
  OAI21X4 U10516 ( .A0(n4860), .A1(n26234), .B0(n4033), .Y(M3_a_11_) );
  AOI21X4 U10517 ( .A0(n25206), .A1(data[43]), .B0(n4655), .Y(n4033) );
  NAND2X1 U10518 ( .A(n3895), .B(n20967), .Y(n4993) );
  INVX8 U10519 ( .A(n25813), .Y(n25206) );
  NAND2X4 U10520 ( .A(n12901), .B(n4948), .Y(n4132) );
  OAI21X1 U10521 ( .A0(n12027), .A1(n12119), .B0(n4040), .Y(n12015) );
  NAND2XL U10522 ( .A(n4968), .B(n4041), .Y(n4040) );
  XOR2X1 U10523 ( .A(n12279), .B(n25884), .Y(n4041) );
  NAND2X1 U10524 ( .A(n5959), .B(n13038), .Y(n4042) );
  NOR2X1 U10525 ( .A(n20668), .B(n4043), .Y(n5959) );
  NAND2XL U10526 ( .A(n12582), .B(n12583), .Y(n4044) );
  NAND2BXL U10527 ( .AN(n12582), .B(n4046), .Y(n4045) );
  XNOR2X1 U10528 ( .A(n12581), .B(n4047), .Y(n12565) );
  XNOR2X1 U10529 ( .A(n12582), .B(n12583), .Y(n4047) );
  INVXL U10530 ( .A(n25915), .Y(n4049) );
  INVX1 U10531 ( .A(n12818), .Y(n4050) );
  NOR2X1 U10532 ( .A(n5959), .B(n13038), .Y(n4053) );
  NAND2X4 U10533 ( .A(n12633), .B(n4054), .Y(n12635) );
  NAND2X1 U10534 ( .A(n12865), .B(n3170), .Y(n4055) );
  AOI21X1 U10535 ( .A0(n12859), .A1(n12863), .B0(n12771), .Y(n12836) );
  OAI22X1 U10536 ( .A0(n11811), .A1(n12597), .B0(n12595), .B1(n4057), .Y(
        n11809) );
  OAI22X1 U10537 ( .A0(n12597), .A1(n4057), .B0(n11674), .B1(n12595), .Y(
        n11732) );
  XNOR2X1 U10538 ( .A(n12594), .B(n12561), .Y(n4057) );
  NAND2X2 U10539 ( .A(n4064), .B(n4062), .Y(n5990) );
  NAND2X2 U10540 ( .A(n17458), .B(n3353), .Y(n4062) );
  NAND2X1 U10541 ( .A(n23751), .B(n3131), .Y(n4064) );
  NAND2X1 U10542 ( .A(n4068), .B(n17933), .Y(n4065) );
  OR2X2 U10543 ( .A(n4068), .B(n17933), .Y(n4066) );
  XOR2X1 U10544 ( .A(n17932), .B(n4067), .Y(n17958) );
  XOR2X1 U10545 ( .A(n4068), .B(n17933), .Y(n4067) );
  NAND2X1 U10546 ( .A(n4069), .B(n5812), .Y(n4068) );
  INVX2 U10547 ( .A(n9739), .Y(n4070) );
  OAI21X1 U10548 ( .A0(n10656), .A1(n10609), .B0(n4072), .Y(n4071) );
  XNOR2X4 U10549 ( .A(n4073), .B(n4940), .Y(n12765) );
  OAI22X1 U10550 ( .A0(n12595), .A1(n12594), .B0(n12597), .B1(n12596), .Y(
        n4075) );
  XOR2X4 U10551 ( .A(n4078), .B(n4678), .Y(n21043) );
  OAI21X4 U10552 ( .A0(n3415), .A1(n12975), .B0(n4079), .Y(n4078) );
  AOI22X1 U10553 ( .A0(n4215), .A1(n24178), .B0(n25502), .B1(n4220), .Y(n4081)
         );
  XOR3X2 U10554 ( .A(n17763), .B(n17764), .C(n17762), .Y(n17798) );
  OAI2BB1X2 U10555 ( .A0N(n17686), .A1N(n4315), .B0(n4082), .Y(n17649) );
  NAND2X1 U10556 ( .A(n17685), .B(n4083), .Y(n4082) );
  NAND2X1 U10557 ( .A(n4316), .B(n4314), .Y(n4083) );
  XOR2X2 U10558 ( .A(n4184), .B(n4182), .Y(n4316) );
  NAND2BX4 U10559 ( .AN(n4085), .B(n4084), .Y(M4_a_17_) );
  NAND2X2 U10560 ( .A(n5015), .B(data[81]), .Y(n4084) );
  OAI22X1 U10561 ( .A0(n17708), .A1(n18625), .B0(n17874), .B1(n18624), .Y(
        n17927) );
  OAI21X2 U10562 ( .A0(n5507), .A1(n18624), .B0(n4086), .Y(n17531) );
  NAND2BX1 U10563 ( .AN(n17507), .B(n3187), .Y(n4086) );
  OAI22X1 U10564 ( .A0(n17693), .A1(n18625), .B0(n18624), .B1(n17708), .Y(
        n17712) );
  NOR2X1 U10565 ( .A(n17517), .B(n17902), .Y(n4088) );
  NOR2X1 U10566 ( .A(n18107), .B(n17581), .Y(n4089) );
  AOI22X2 U10567 ( .A0(n25590), .A1(n4220), .B0(n4215), .B1(n23479), .Y(n24129) );
  XOR2X2 U10568 ( .A(n16973), .B(n4098), .Y(n16995) );
  XOR2X1 U10569 ( .A(n16974), .B(n4099), .Y(n4098) );
  OAI22X1 U10570 ( .A0(n16941), .A1(n16940), .B0(n16939), .B1(n3203), .Y(n4099) );
  OAI21X2 U10571 ( .A0(n17316), .A1(n17314), .B0(n17317), .Y(n17312) );
  AOI21X1 U10572 ( .A0(n17363), .A1(n5667), .B0(n17362), .Y(n17364) );
  INVX1 U10573 ( .A(n3085), .Y(n4105) );
  AOI21X4 U10574 ( .A0(n5666), .A1(n5667), .B0(n4107), .Y(n4106) );
  OAI22XL U10575 ( .A0(n16941), .A1(n16342), .B0(n16939), .B1(n4109), .Y(
        n16366) );
  NOR2X1 U10576 ( .A(n16941), .B(n4109), .Y(n4108) );
  XOR2X1 U10577 ( .A(n5430), .B(n16873), .Y(n4109) );
  NAND2XL U10578 ( .A(n16448), .B(n16449), .Y(n4110) );
  OR2X2 U10579 ( .A(n16448), .B(n16449), .Y(n4111) );
  XNOR2X2 U10580 ( .A(n16447), .B(n4112), .Y(n16452) );
  AOI21X4 U10581 ( .A0(n10125), .A1(n10198), .B0(n4114), .Y(n10126) );
  OAI21X2 U10582 ( .A0(n10201), .A1(n10206), .B0(n10202), .Y(n4114) );
  XOR2X4 U10583 ( .A(n4115), .B(n3008), .Y(n10122) );
  NOR2X4 U10584 ( .A(n10201), .B(n10200), .Y(n10125) );
  AND2X4 U10585 ( .A(n4116), .B(n5062), .Y(n23643) );
  AOI21X4 U10586 ( .A0(n10191), .A1(n5235), .B0(n4117), .Y(n5234) );
  OAI21X4 U10587 ( .A0(n10230), .A1(n10237), .B0(n10238), .Y(n4117) );
  NOR2X4 U10588 ( .A(n10195), .B(n10237), .Y(n5235) );
  NOR2X4 U10589 ( .A(n10142), .B(n10143), .Y(n10237) );
  OAI21X4 U10590 ( .A0(n10186), .A1(n10223), .B0(n10187), .Y(n10191) );
  NAND2X2 U10591 ( .A(n10139), .B(n10138), .Y(n10187) );
  NAND2X2 U10592 ( .A(n10137), .B(n10136), .Y(n10223) );
  NOR2X4 U10593 ( .A(n10139), .B(n10138), .Y(n10186) );
  OAI21X4 U10594 ( .A0(n4120), .A1(n4119), .B0(n4118), .Y(n9556) );
  XNOR3X4 U10595 ( .A(n9509), .B(n9508), .C(n4120), .Y(n9490) );
  XNOR3X2 U10596 ( .A(n9523), .B(n9521), .C(n9522), .Y(n4120) );
  NAND2XL U10597 ( .A(n3132), .B(n4121), .Y(n5315) );
  INVX1 U10598 ( .A(n19048), .Y(n4121) );
  INVX1 U10599 ( .A(n23750), .Y(n4122) );
  NAND2X4 U10600 ( .A(n5343), .B(n9838), .Y(n9551) );
  XNOR2X4 U10601 ( .A(M2_a_6_), .B(M2_a_5_), .Y(n9838) );
  NAND3BX4 U10602 ( .AN(n5348), .B(n9062), .C(n4124), .Y(M2_a_5_) );
  OAI22XL U10603 ( .A0(n3102), .A1(n4126), .B0(n16165), .B1(n16332), .Y(n16161) );
  INVX1 U10604 ( .A(n4129), .Y(n4127) );
  INVX1 U10605 ( .A(n12432), .Y(n4133) );
  INVXL U10606 ( .A(n3183), .Y(n4134) );
  OAI21XL U10607 ( .A0(n16172), .A1(n16173), .B0(n16171), .Y(n4136) );
  NOR2X2 U10608 ( .A(n10057), .B(n10058), .Y(n4141) );
  NAND2X1 U10609 ( .A(n10056), .B(n10055), .Y(n4140) );
  OAI2BB1X2 U10610 ( .A0N(n13979), .A1N(n4146), .B0(n4144), .Y(n14005) );
  NAND2X1 U10611 ( .A(n13978), .B(n4145), .Y(n4144) );
  OR2XL U10612 ( .A(n13979), .B(n4146), .Y(n4145) );
  NAND2X1 U10613 ( .A(n4874), .B(n4147), .Y(n4146) );
  OAI21XL U10614 ( .A0(n13928), .A1(n13927), .B0(n13926), .Y(n4147) );
  OAI21X1 U10615 ( .A0(n13917), .A1(n14268), .B0(n4148), .Y(n13927) );
  OR2X2 U10616 ( .A(n13900), .B(n14282), .Y(n4148) );
  OAI2BB1X2 U10617 ( .A0N(n17236), .A1N(n17304), .B0(n3158), .Y(n4149) );
  NAND2X1 U10618 ( .A(n17304), .B(n17297), .Y(n4151) );
  NAND2X1 U10619 ( .A(n3081), .B(n4155), .Y(n4300) );
  NAND3X1 U10620 ( .A(n3081), .B(n4155), .C(n25786), .Y(n4302) );
  AOI22X1 U10621 ( .A0(n3081), .A1(n23879), .B0(n4267), .B1(n4155), .Y(n24145)
         );
  OAI21XL U10622 ( .A0(n16000), .A1(n5808), .B0(n15999), .Y(n5807) );
  NAND2XL U10623 ( .A(n4165), .B(n5760), .Y(n4156) );
  NOR2XL U10624 ( .A(n16011), .B(n16942), .Y(n4157) );
  NAND2BX4 U10625 ( .AN(n20677), .B(n4158), .Y(n5157) );
  NOR2X2 U10626 ( .A(n17230), .B(n17231), .Y(n17249) );
  NOR2X2 U10627 ( .A(n16851), .B(n16850), .Y(n17230) );
  CLKINVX3 U10628 ( .A(n17465), .Y(n20919) );
  XOR2X4 U10629 ( .A(n4161), .B(n17386), .Y(n17465) );
  XOR2X2 U10630 ( .A(n16967), .B(n3176), .Y(n4162) );
  XNOR3X2 U10631 ( .A(n4166), .B(n16964), .C(n6013), .Y(n5725) );
  OAI21X2 U10632 ( .A0(n16942), .A1(n15968), .B0(n4163), .Y(n16964) );
  XOR2X1 U10633 ( .A(n6162), .B(n18468), .Y(n17582) );
  NAND2X1 U10634 ( .A(n3136), .B(n21048), .Y(n4167) );
  OAI22X1 U10635 ( .A0(n4169), .A1(n16475), .B0(n16108), .B1(n16638), .Y(
        n16425) );
  INVX1 U10636 ( .A(n4170), .Y(n18895) );
  NOR2X2 U10637 ( .A(n4170), .B(n4207), .Y(n18422) );
  XOR2X1 U10638 ( .A(M4_a_17_), .B(n4206), .Y(n18444) );
  XOR2X1 U10639 ( .A(n18638), .B(n4206), .Y(n18481) );
  XOR2X1 U10640 ( .A(n18500), .B(n4206), .Y(n17783) );
  XNOR2X1 U10641 ( .A(n16614), .B(n18673), .Y(n15958) );
  XOR2XL U10642 ( .A(n18468), .B(n4206), .Y(n18434) );
  XOR2X1 U10643 ( .A(n18118), .B(n4206), .Y(n17504) );
  XOR2X1 U10644 ( .A(n18453), .B(n4206), .Y(n18540) );
  XOR2X1 U10645 ( .A(n18658), .B(n18673), .Y(n4200) );
  XNOR2XL U10646 ( .A(n18150), .B(M3_mult_x_15_b_20_), .Y(n17520) );
  XNOR2X1 U10647 ( .A(n5729), .B(n4206), .Y(n4177) );
  XOR2X2 U10648 ( .A(n6081), .B(n4171), .Y(n4509) );
  NAND2X1 U10649 ( .A(n20659), .B(n25796), .Y(n4172) );
  XOR2X1 U10650 ( .A(n9366), .B(n9367), .Y(n4176) );
  NAND2X2 U10651 ( .A(n4657), .B(n4178), .Y(n9335) );
  OAI21XL U10652 ( .A0(n9279), .A1(n4321), .B0(n9278), .Y(n4178) );
  OAI21X2 U10653 ( .A0(n10496), .A1(n9217), .B0(n4339), .Y(n4321) );
  NAND2X1 U10654 ( .A(n4179), .B(n5506), .Y(n18325) );
  NAND3X2 U10655 ( .A(n4181), .B(n5473), .C(n4180), .Y(n25379) );
  NAND2X1 U10656 ( .A(n5888), .B(n5771), .Y(n4180) );
  NAND2BX2 U10657 ( .AN(n5888), .B(n5009), .Y(n4181) );
  INVX1 U10658 ( .A(n17592), .Y(n4182) );
  XOR2X1 U10659 ( .A(n17593), .B(n17594), .Y(n4184) );
  NAND2X1 U10660 ( .A(n4185), .B(n5446), .Y(n23732) );
  NAND2XL U10661 ( .A(n4185), .B(n23734), .Y(n23511) );
  NOR2X4 U10662 ( .A(n4203), .B(n3146), .Y(n4185) );
  OAI21XL U10663 ( .A0(n17604), .A1(n17962), .B0(n4186), .Y(n17680) );
  OAI21X1 U10664 ( .A0(n17715), .A1(n18177), .B0(n4187), .Y(n17868) );
  NOR2BXL U10665 ( .AN(n18428), .B(n4189), .Y(M4_U3_U1_enc_tree_1__1__20_) );
  AOI21XL U10666 ( .A0(n18110), .A1(n4189), .B0(n4196), .Y(
        M4_U3_U1_enc_tree_0__1__22_) );
  NAND3BX4 U10667 ( .AN(n5031), .B(n4398), .C(n4660), .Y(n4189) );
  NAND2X2 U10668 ( .A(n4192), .B(n4830), .Y(n10114) );
  OAI21XL U10669 ( .A0(n9684), .A1(n9686), .B0(n9685), .Y(n4192) );
  NAND2X2 U10670 ( .A(n6067), .B(n6068), .Y(n9684) );
  OAI22XL U10671 ( .A0(n10496), .A1(n9603), .B0(n9504), .B1(n9652), .Y(n9633)
         );
  XOR2X1 U10672 ( .A(n6076), .B(M2_a_17_), .Y(n9652) );
  OR2X2 U10673 ( .A(n18363), .B(n18364), .Y(n4194) );
  XOR3X2 U10674 ( .A(n18362), .B(n18363), .C(n18364), .Y(n18382) );
  XOR2X2 U10675 ( .A(M4_a_7_), .B(n4196), .Y(n4195) );
  XOR2X1 U10676 ( .A(M4_a_9_), .B(n4196), .Y(n4519) );
  NOR2BXL U10677 ( .AN(n4197), .B(n18830), .Y(n24251) );
  NAND2BXL U10678 ( .AN(n5475), .B(n4197), .Y(n24253) );
  AOI21X2 U10679 ( .A0(n4198), .A1(n20655), .B0(n20653), .Y(n5439) );
  XNOR2X4 U10680 ( .A(n4375), .B(n4699), .Y(n5437) );
  NAND2X1 U10681 ( .A(n18962), .B(n18966), .Y(n18703) );
  OAI22X1 U10682 ( .A0(n18659), .A1(n18609), .B0(n17832), .B1(n4200), .Y(
        n18619) );
  NAND2X2 U10683 ( .A(n18411), .B(n18410), .Y(n18899) );
  NOR2X4 U10684 ( .A(n18412), .B(n18413), .Y(n18890) );
  OAI21X4 U10685 ( .A0(n19014), .A1(n18853), .B0(n18852), .Y(n4202) );
  NOR2X4 U10686 ( .A(n4404), .B(n23476), .Y(n23527) );
  NAND2BX1 U10687 ( .AN(n17743), .B(n3104), .Y(n4204) );
  OAI22X1 U10688 ( .A0(n17621), .A1(n18111), .B0(n18504), .B1(n4205), .Y(
        n17729) );
  XOR2X1 U10689 ( .A(n4206), .B(n18503), .Y(n4205) );
  OAI21X1 U10690 ( .A0(n18866), .A1(n4207), .B0(n18420), .Y(n18421) );
  NAND2X2 U10691 ( .A(n18865), .B(n18419), .Y(n4207) );
  OAI21X1 U10692 ( .A0(n17730), .A1(n4209), .B0(n4208), .Y(n5796) );
  NAND2XL U10693 ( .A(n5797), .B(n17730), .Y(n4208) );
  NOR2X1 U10694 ( .A(n5798), .B(n4211), .Y(n5797) );
  NOR2X1 U10695 ( .A(n4211), .B(n5798), .Y(n4209) );
  OAI22X1 U10696 ( .A0(n17619), .A1(n18624), .B0(n17748), .B1(n18625), .Y(
        n17730) );
  CLKINVX8 U10697 ( .A(n18106), .Y(n18118) );
  INVX8 U10698 ( .A(n18603), .Y(n18604) );
  NOR2X1 U10699 ( .A(n17735), .B(n17902), .Y(n4211) );
  XOR2X1 U10700 ( .A(n18106), .B(n3202), .Y(n17735) );
  XOR2X1 U10701 ( .A(n18603), .B(n12561), .Y(n17748) );
  NOR2X4 U10702 ( .A(n4511), .B(n4510), .Y(n4210) );
  AOI22X2 U10703 ( .A0(n4215), .A1(n25528), .B0(n4220), .B1(n25552), .Y(n24147) );
  NAND2X1 U10704 ( .A(n23734), .B(n23528), .Y(n4214) );
  NAND2X1 U10705 ( .A(n3014), .B(n4222), .Y(n4217) );
  XOR2X2 U10706 ( .A(n23520), .B(n23519), .Y(n24179) );
  NOR2X4 U10707 ( .A(n4225), .B(n4224), .Y(n18658) );
  NOR2X1 U10708 ( .A(n25813), .B(n26265), .Y(n4226) );
  INVX1 U10709 ( .A(n12420), .Y(n4228) );
  NAND2XL U10710 ( .A(n12405), .B(n12406), .Y(n4230) );
  NAND2BX1 U10711 ( .AN(n12407), .B(n4234), .Y(n4231) );
  OAI21XL U10712 ( .A0(n12404), .A1(n12403), .B0(n4234), .Y(n4233) );
  AOI21X1 U10713 ( .A0(n12382), .A1(n12383), .B0(n12381), .Y(n4235) );
  OAI22XL U10714 ( .A0(n12186), .A1(n12338), .B0(n12340), .B1(n4238), .Y(
        n12206) );
  XOR2X1 U10715 ( .A(n16884), .B(n4239), .Y(n4238) );
  INVXL U10716 ( .A(n2980), .Y(n4239) );
  AOI22XL U10717 ( .A0(n23795), .A1(n25294), .B0(temp1[1]), .B1(n2983), .Y(
        n23441) );
  NAND2X4 U10718 ( .A(n4343), .B(n17902), .Y(n18107) );
  NAND2X2 U10719 ( .A(n4242), .B(n5892), .Y(M4_a_6_) );
  AOI22X1 U10720 ( .A0(n4875), .A1(data[70]), .B0(in_valid_t), .B1(w2[38]), 
        .Y(n4242) );
  AOI22X1 U10721 ( .A0(n5770), .A1(data[69]), .B0(in_valid_t), .B1(w2[37]), 
        .Y(n4243) );
  NOR2BX1 U10722 ( .AN(n23489), .B(n23736), .Y(n23737) );
  NOR2X2 U10723 ( .A(n4245), .B(n3078), .Y(n5012) );
  NOR2X1 U10724 ( .A(n4245), .B(n5526), .Y(n5525) );
  OAI21XL U10725 ( .A0(n18558), .A1(n18559), .B0(n18557), .Y(n4246) );
  XNOR3X2 U10726 ( .A(n18559), .B(n18558), .C(n4247), .Y(n18586) );
  NOR2X1 U10727 ( .A(n4248), .B(n18942), .Y(n18960) );
  NOR2X1 U10728 ( .A(n4248), .B(n18983), .Y(n18999) );
  OAI21X1 U10729 ( .A0(n19014), .A1(n4248), .B0(n18984), .Y(n18943) );
  AND2X4 U10730 ( .A(n18694), .B(n18846), .Y(n19007) );
  OAI22X1 U10731 ( .A0(n17825), .A1(n18624), .B0(n18625), .B1(n4249), .Y(
        n18534) );
  OAI22X1 U10732 ( .A0(n18499), .A1(n18625), .B0(n18624), .B1(n4249), .Y(
        n18537) );
  OAI22X1 U10733 ( .A0(n10517), .A1(n9599), .B0(n10533), .B1(n6075), .Y(n9611)
         );
  XOR2X1 U10734 ( .A(n10494), .B(n6076), .Y(n6075) );
  NOR2X2 U10735 ( .A(n5499), .B(n14662), .Y(n23480) );
  OAI2BB1X4 U10736 ( .A0N(n4939), .A1N(n4263), .B0(n4253), .Y(n5499) );
  XOR2X1 U10737 ( .A(n25864), .B(n4254), .Y(n13430) );
  OAI21X4 U10738 ( .A0(n3115), .A1(n25916), .B0(n11540), .Y(n25864) );
  OAI21X1 U10739 ( .A0(n24115), .A1(n5770), .B0(n24114), .Y(n4255) );
  NOR2X1 U10740 ( .A(n5917), .B(n4257), .Y(n4256) );
  NAND3XL U10741 ( .A(n4258), .B(n14398), .C(n3152), .Y(n4484) );
  AOI21XL U10742 ( .A0(n4258), .A1(n14398), .B0(n14397), .Y(n14402) );
  NAND2X2 U10743 ( .A(n4267), .B(n23592), .Y(n4259) );
  OAI21XL U10744 ( .A0(n13309), .A1(n13310), .B0(n13308), .Y(n4260) );
  XOR3X2 U10745 ( .A(n13310), .B(n13308), .C(n13309), .Y(n13250) );
  NOR2X2 U10746 ( .A(n13998), .B(n13999), .Y(n14585) );
  NAND2X1 U10747 ( .A(n24655), .B(n4579), .Y(n4978) );
  NAND2X1 U10748 ( .A(n4267), .B(n23631), .Y(n4264) );
  XOR2X1 U10749 ( .A(M1_b_8_), .B(n14043), .Y(n13041) );
  INVX1 U10750 ( .A(n6210), .Y(n14043) );
  AOI21X4 U10751 ( .A0(n25233), .A1(learning_rate[9]), .B0(n4265), .Y(n6210)
         );
  NAND2X2 U10752 ( .A(n13040), .B(n5166), .Y(n4265) );
  NAND2X2 U10753 ( .A(n4479), .B(n4266), .Y(M1_b_8_) );
  NAND2X1 U10754 ( .A(n25233), .B(learning_rate[8]), .Y(n4266) );
  NAND3X1 U10755 ( .A(n23441), .B(n23440), .C(n4268), .Y(n2553) );
  OR2X2 U10756 ( .A(n5085), .B(n4583), .Y(n4268) );
  AOI22X2 U10757 ( .A0(n23592), .A1(n3081), .B0(n4267), .B1(n23483), .Y(n5085)
         );
  AOI21X4 U10758 ( .A0(n14551), .A1(n14556), .B0(n4269), .Y(n14520) );
  NAND2X1 U10759 ( .A(n14315), .B(n14316), .Y(n14555) );
  NAND2X4 U10760 ( .A(n4271), .B(n4270), .Y(n14556) );
  CLKINVX3 U10761 ( .A(n14316), .Y(n4270) );
  XOR2X4 U10762 ( .A(n5489), .B(M1_b_12_), .Y(n14120) );
  NAND2X4 U10763 ( .A(n4273), .B(n4272), .Y(M1_b_12_) );
  NAND2XL U10764 ( .A(n4275), .B(n14083), .Y(n4274) );
  XOR2X1 U10765 ( .A(n14084), .B(n4277), .Y(n14104) );
  NOR2X1 U10766 ( .A(n4280), .B(n4279), .Y(n4278) );
  NOR2X1 U10767 ( .A(n14157), .B(n14070), .Y(n4279) );
  NOR2XL U10768 ( .A(n5510), .B(n14120), .Y(n4280) );
  NAND2X1 U10769 ( .A(n4281), .B(n3083), .Y(n20689) );
  NOR2X1 U10770 ( .A(n20687), .B(n3134), .Y(n4281) );
  NAND3X1 U10771 ( .A(n6109), .B(n6108), .C(n4282), .Y(n2532) );
  NOR2X1 U10772 ( .A(n13343), .B(n13342), .Y(n13346) );
  NAND2X2 U10773 ( .A(n5274), .B(n4284), .Y(n23431) );
  INVXL U10774 ( .A(n4284), .Y(n4294) );
  NAND2XL U10775 ( .A(n20973), .B(n4284), .Y(n23445) );
  OAI21X4 U10776 ( .A0(n3103), .A1(n4287), .B0(n4285), .Y(M1_b_3_) );
  NOR2BX4 U10777 ( .AN(n5089), .B(n4286), .Y(n4285) );
  AND3X4 U10778 ( .A(n13356), .B(n4290), .C(n4289), .Y(n4288) );
  NAND2X1 U10779 ( .A(in_valid_d), .B(w1[145]), .Y(n4289) );
  NAND2X1 U10780 ( .A(n4566), .B(learning_rate[17]), .Y(n4290) );
  CLKINVX8 U10781 ( .A(n5157), .Y(n23744) );
  INVX1 U10782 ( .A(n20328), .Y(n4292) );
  NOR2X1 U10783 ( .A(n5157), .B(n4294), .Y(n4293) );
  NAND2XL U10784 ( .A(n5211), .B(n23568), .Y(n4295) );
  NOR2BX1 U10785 ( .AN(n20981), .B(n5157), .Y(n4296) );
  AOI21X1 U10786 ( .A0(n14647), .A1(n14511), .B0(n14510), .Y(n14512) );
  OAI21X2 U10787 ( .A0(n14533), .A1(n14503), .B0(n14502), .Y(n14647) );
  AOI21X4 U10788 ( .A0(n14322), .A1(n14552), .B0(n4297), .Y(n14533) );
  OAI21X4 U10789 ( .A0(n14520), .A1(n5494), .B0(n5392), .Y(n4297) );
  OAI21X2 U10790 ( .A0(n14573), .A1(n14591), .B0(n14574), .Y(n14552) );
  NOR2X4 U10791 ( .A(n14521), .B(n5494), .Y(n14322) );
  OAI22XL U10792 ( .A0(n14023), .A1(n14249), .B0(n14250), .B1(n4298), .Y(
        n14050) );
  NAND2X1 U10793 ( .A(n4300), .B(n4299), .Y(n24555) );
  NAND2X1 U10794 ( .A(n4267), .B(n23569), .Y(n4299) );
  NAND2X1 U10795 ( .A(n4302), .B(n4301), .Y(n24144) );
  NAND3X1 U10796 ( .A(n4267), .B(n23569), .C(n25786), .Y(n4301) );
  XOR3X2 U10797 ( .A(n9283), .B(n9284), .C(n9285), .Y(n9373) );
  OAI21X1 U10798 ( .A0(n9983), .A1(n4303), .B0(n4312), .Y(n4311) );
  OAI22X1 U10799 ( .A0(n9983), .A1(n9253), .B0(n9906), .B1(n4303), .Y(n9259)
         );
  NAND2XL U10800 ( .A(n20610), .B(n4305), .Y(n17486) );
  NAND2XL U10801 ( .A(n9246), .B(n4311), .Y(n4307) );
  XNOR3X2 U10802 ( .A(n17686), .B(n4316), .C(n17685), .Y(n17687) );
  INVXL U10803 ( .A(n17596), .Y(n4317) );
  NAND2X4 U10804 ( .A(n4318), .B(n13427), .Y(n14282) );
  CLKINVX3 U10805 ( .A(n13428), .Y(n4318) );
  XNOR2X1 U10806 ( .A(n12667), .B(n12668), .Y(n5041) );
  XOR2X1 U10807 ( .A(n3202), .B(M3_U3_U1_or2_inv_0__18_), .Y(n4890) );
  NAND3XL U10808 ( .A(n20666), .B(n4320), .C(n23706), .Y(n23708) );
  NAND2X1 U10809 ( .A(n20666), .B(n4320), .Y(n20661) );
  AND2X2 U10810 ( .A(n20665), .B(n14689), .Y(n4320) );
  XOR3X2 U10811 ( .A(n9279), .B(n4321), .C(n9278), .Y(n9287) );
  NOR2XL U10812 ( .A(n10341), .B(n10311), .Y(M2_U4_U1_or2_tree_0__1__20_) );
  INVX4 U10813 ( .A(M2_U4_U1_or2_inv_0__22_), .Y(n10311) );
  AND2X2 U10814 ( .A(n3895), .B(n21032), .Y(n4967) );
  OAI21XL U10815 ( .A0(n9368), .A1(n9367), .B0(n9366), .Y(n4323) );
  NAND2BX2 U10816 ( .AN(n10054), .B(n3091), .Y(n4325) );
  NOR2X2 U10817 ( .A(n20944), .B(n4690), .Y(n4326) );
  NOR2X2 U10818 ( .A(n6071), .B(n10198), .Y(n4327) );
  NAND2XL U10819 ( .A(n4331), .B(n17484), .Y(n23491) );
  XOR2X1 U10820 ( .A(n9715), .B(n9717), .Y(n5142) );
  XOR2X1 U10821 ( .A(n9892), .B(n6076), .Y(n4334) );
  OAI21X4 U10822 ( .A0(n18919), .A1(n4507), .B0(n18920), .Y(n18904) );
  OR2X2 U10823 ( .A(n17704), .B(n17703), .Y(n4337) );
  OAI22X1 U10824 ( .A0(n18652), .A1(n4338), .B0(n17872), .B1(n17529), .Y(
        n17587) );
  OAI22X1 U10825 ( .A0(n18652), .A1(n17674), .B0(n17872), .B1(n4338), .Y(
        n17700) );
  XOR2X1 U10826 ( .A(n18638), .B(n3114), .Y(n4338) );
  INVXL U10827 ( .A(n9287), .Y(n4817) );
  BUFX3 U10828 ( .A(n19043), .Y(n4342) );
  NOR2X1 U10829 ( .A(n19043), .B(n3111), .Y(n5269) );
  XNOR2X4 U10830 ( .A(n10633), .B(n10632), .Y(n17485) );
  NAND2X1 U10831 ( .A(n20685), .B(n4344), .Y(n20686) );
  NAND2XL U10832 ( .A(n19072), .B(n3066), .Y(n4346) );
  NAND2X1 U10833 ( .A(n3128), .B(n19075), .Y(n4348) );
  INVX1 U10834 ( .A(n9740), .Y(n4349) );
  XOR3X2 U10835 ( .A(n9740), .B(n9739), .C(n9738), .Y(n9765) );
  NAND2X2 U10836 ( .A(n6071), .B(n3151), .Y(n4350) );
  AOI21X1 U10837 ( .A0(n10198), .A1(n3151), .B0(n4352), .Y(n4351) );
  NAND3X1 U10838 ( .A(n5741), .B(n10718), .C(n6074), .Y(n19054) );
  OAI21X4 U10839 ( .A0(n19053), .A1(n20947), .B0(n19054), .Y(n23738) );
  CLKINVX3 U10840 ( .A(n10718), .Y(n5174) );
  NAND2XL U10841 ( .A(n2976), .B(n4357), .Y(n4354) );
  XOR2X1 U10842 ( .A(n2976), .B(n4357), .Y(n4356) );
  OAI2BB1X2 U10843 ( .A0N(n5183), .A1N(n6164), .B0(n10429), .Y(n4359) );
  OAI2BB1X2 U10844 ( .A0N(n3122), .A1N(n24606), .B0(n24599), .Y(n24600) );
  NAND2X2 U10845 ( .A(n4362), .B(n4361), .Y(n24606) );
  NAND2X1 U10846 ( .A(n23926), .B(n3128), .Y(n4361) );
  NAND2X1 U10847 ( .A(n23925), .B(n19104), .Y(n4362) );
  XOR2X4 U10848 ( .A(n4367), .B(n4624), .Y(n21039) );
  OAI21X4 U10849 ( .A0(n3415), .A1(n12847), .B0(n12846), .Y(n4368) );
  NAND2X4 U10850 ( .A(n4369), .B(n20648), .Y(n24386) );
  NOR2X1 U10851 ( .A(n4369), .B(n20645), .Y(n5352) );
  OAI21XL U10852 ( .A0(n20798), .A1(n4369), .B0(n24380), .Y(n20804) );
  OAI21XL U10853 ( .A0(n20779), .A1(n4369), .B0(n24380), .Y(n20783) );
  OAI21XL U10854 ( .A0(n23659), .A1(n4369), .B0(n24380), .Y(n23666) );
  OAI21XL U10855 ( .A0(n23774), .A1(n4369), .B0(n24380), .Y(n23780) );
  OAI21XL U10856 ( .A0(n24381), .A1(n4369), .B0(n24380), .Y(n24388) );
  OAI21XL U10857 ( .A0(n24267), .A1(n4369), .B0(n24380), .Y(n24273) );
  NAND2X4 U10858 ( .A(n4369), .B(n20644), .Y(n24380) );
  NAND2X4 U10859 ( .A(n4463), .B(n5173), .Y(n4369) );
  NAND3BX2 U10860 ( .AN(n6106), .B(n4645), .C(n20353), .Y(n25331) );
  XNOR3X2 U10861 ( .A(n4373), .B(n4372), .C(n17770), .Y(n17804) );
  INVXL U10862 ( .A(n17771), .Y(n4372) );
  XOR2X1 U10863 ( .A(n5886), .B(n17740), .Y(n4373) );
  NAND2X4 U10864 ( .A(n23561), .B(n4374), .Y(n23734) );
  OAI21X4 U10865 ( .A0(n19014), .A1(n18719), .B0(n18718), .Y(n4375) );
  NAND2X1 U10866 ( .A(n4376), .B(n12218), .Y(n12420) );
  AOI21X1 U10867 ( .A0(n12418), .A1(n4376), .B0(n12417), .Y(n12419) );
  NOR2X1 U10868 ( .A(n3014), .B(n5771), .Y(n5009) );
  NAND2X1 U10869 ( .A(n3014), .B(n5771), .Y(n5473) );
  XOR2X4 U10870 ( .A(n4377), .B(n4684), .Y(n13024) );
  OAI21X1 U10871 ( .A0(n12598), .A1(n4381), .B0(n6009), .Y(n12185) );
  OAI21XL U10872 ( .A0(n12342), .A1(n4381), .B0(n4384), .Y(n12390) );
  XOR2X1 U10873 ( .A(n3204), .B(n3114), .Y(n4381) );
  XOR2X2 U10874 ( .A(n5966), .B(n13025), .Y(n4382) );
  OAI21XL U10875 ( .A0(n12341), .A1(n12598), .B0(n4383), .Y(n12334) );
  NAND2XL U10876 ( .A(n4385), .B(n3186), .Y(n4383) );
  NAND2XL U10877 ( .A(n4385), .B(n3709), .Y(n4384) );
  XOR2X1 U10878 ( .A(n12279), .B(n3204), .Y(n4385) );
  NAND2XL U10879 ( .A(n12404), .B(n12403), .Y(n12407) );
  NAND2X1 U10880 ( .A(n4387), .B(n4386), .Y(n12386) );
  NAND2XL U10881 ( .A(n12395), .B(n12396), .Y(n4386) );
  NAND2X1 U10882 ( .A(n4388), .B(n12394), .Y(n4387) );
  OR2X2 U10883 ( .A(n12395), .B(n12396), .Y(n4388) );
  XOR2X1 U10884 ( .A(n12395), .B(n4389), .Y(n12397) );
  XOR2X1 U10885 ( .A(n12396), .B(n12394), .Y(n4389) );
  NAND3X1 U10886 ( .A(n3894), .B(n5978), .C(n17456), .Y(n5402) );
  NAND2XL U10887 ( .A(n17940), .B(n4394), .Y(n4390) );
  XOR2X1 U10888 ( .A(n17940), .B(n4394), .Y(n4393) );
  NAND2X4 U10889 ( .A(n18501), .B(n4396), .Y(n18083) );
  NAND2X1 U10890 ( .A(n5032), .B(data[73]), .Y(n4397) );
  OAI2BB1X2 U10891 ( .A0N(n18009), .A1N(n4401), .B0(n4399), .Y(n17987) );
  NAND2X1 U10892 ( .A(n4400), .B(n18010), .Y(n4399) );
  NAND2X1 U10893 ( .A(n4403), .B(n4402), .Y(n4401) );
  INVXL U10894 ( .A(n18010), .Y(n4402) );
  XNOR3X2 U10895 ( .A(n18010), .B(n4403), .C(n18009), .Y(n18011) );
  OAI21X1 U10896 ( .A0(n18925), .A1(n18913), .B0(n18912), .Y(n4406) );
  XOR3X2 U10897 ( .A(n18361), .B(n18360), .C(n18359), .Y(n18388) );
  NAND2XL U10898 ( .A(n4422), .B(n4423), .Y(n4421) );
  NOR2X1 U10899 ( .A(n11829), .B(n12718), .Y(n4424) );
  NOR2X1 U10900 ( .A(n11843), .B(n12717), .Y(n4425) );
  XOR2X1 U10901 ( .A(n4430), .B(n11718), .Y(n11863) );
  OAI22X2 U10902 ( .A0(n12759), .A1(n5976), .B0(n12760), .B1(n11917), .Y(
        n11922) );
  XNOR2X1 U10903 ( .A(n12758), .B(M3_mult_x_15_b_9_), .Y(n11917) );
  NOR2X1 U10904 ( .A(n25796), .B(n26243), .Y(n4432) );
  NAND2X4 U10905 ( .A(n11626), .B(n12222), .Y(n12352) );
  NAND2XL U10906 ( .A(n4440), .B(n12542), .Y(n4435) );
  XOR2X1 U10907 ( .A(n12541), .B(n4439), .Y(n12536) );
  OAI22X1 U10908 ( .A0(n12535), .A1(n12518), .B0(n12995), .B1(n12701), .Y(
        n4440) );
  NOR2XL U10909 ( .A(n20990), .B(n4442), .Y(n20987) );
  NAND2XL U10910 ( .A(n11730), .B(n4448), .Y(n4444) );
  INVXL U10911 ( .A(n4448), .Y(n4446) );
  XOR2X2 U10912 ( .A(n11729), .B(n4447), .Y(n11806) );
  XOR2X1 U10913 ( .A(n11730), .B(n4448), .Y(n4447) );
  OAI22X1 U10914 ( .A0(n11662), .A1(n12760), .B0(n12759), .B1(n11728), .Y(
        n4448) );
  NOR2X1 U10915 ( .A(n15759), .B(n15755), .Y(n15695) );
  NAND2X1 U10916 ( .A(n15757), .B(n23955), .Y(n15759) );
  NAND3XL U10917 ( .A(n15835), .B(n15836), .C(n15772), .Y(n4453) );
  AOI2BB1XL U10918 ( .A0N(n15706), .A1N(n15823), .B0(n4454), .Y(n15707) );
  INVXL U10919 ( .A(n15825), .Y(n4454) );
  NAND2X1 U10920 ( .A(n25269), .B(n23966), .Y(n15746) );
  AOI2BB1X4 U10921 ( .A0N(n4455), .A1N(n25268), .B0(n15782), .Y(n25269) );
  NAND2XL U10922 ( .A(n15277), .B(n3016), .Y(n15312) );
  NOR2XL U10923 ( .A(n4460), .B(n15920), .Y(n15714) );
  OAI21XL U10924 ( .A0(n4462), .A1(n15860), .B0(n15713), .Y(n4461) );
  NOR2XL U10925 ( .A(n15712), .B(n15861), .Y(n4462) );
  NAND3X2 U10926 ( .A(n5232), .B(n5231), .C(n5233), .Y(n4463) );
  INVXL U10927 ( .A(n11531), .Y(n4465) );
  NAND2X4 U10928 ( .A(n4467), .B(n14905), .Y(n15008) );
  XOR2X2 U10929 ( .A(n10066), .B(n10067), .Y(n4468) );
  NAND2X1 U10930 ( .A(n5032), .B(n4732), .Y(n4469) );
  NAND2X2 U10931 ( .A(n5153), .B(n4470), .Y(n4471) );
  NAND2X2 U10932 ( .A(n23568), .B(n3081), .Y(n4470) );
  NAND2XL U10933 ( .A(n3065), .B(n4471), .Y(n5406) );
  AND2X2 U10934 ( .A(n4471), .B(n3060), .Y(n4672) );
  AOI21XL U10935 ( .A0(n25754), .A1(n4471), .B0(n24130), .Y(n2305) );
  NAND2X2 U10936 ( .A(n4476), .B(n14692), .Y(n4475) );
  NOR2X1 U10937 ( .A(n13346), .B(n4477), .Y(n13339) );
  CLKINVX2 U10938 ( .A(n14045), .Y(n13051) );
  XNOR2X1 U10939 ( .A(M1_b_8_), .B(n4807), .Y(n14045) );
  NAND2X4 U10940 ( .A(n5295), .B(n4478), .Y(n4807) );
  NAND2X1 U10941 ( .A(n4579), .B(w1[136]), .Y(n4480) );
  XOR2X2 U10942 ( .A(M1_b_10_), .B(n6210), .Y(n14081) );
  INVXL U10943 ( .A(n14400), .Y(n4483) );
  AOI21XL U10944 ( .A0(n4485), .A1(M3_mult_x_15_b_6_), .B0(n11499), .Y(
        M3_U4_U1_enc_tree_0__1__26_) );
  INVXL U10945 ( .A(n2974), .Y(n4485) );
  NAND2BXL U10946 ( .AN(n12176), .B(n6004), .Y(n4486) );
  OAI22X1 U10947 ( .A0(n4490), .A1(n4489), .B0(n4488), .B1(n4487), .Y(n17670)
         );
  NOR2X1 U10948 ( .A(n17586), .B(n17832), .Y(n4491) );
  XNOR3X2 U10949 ( .A(n4496), .B(n13501), .C(n13500), .Y(n13505) );
  INVX1 U10950 ( .A(n13502), .Y(n4496) );
  NAND2X1 U10951 ( .A(n24048), .B(n25184), .Y(n4497) );
  NAND2X1 U10952 ( .A(n3005), .B(n25185), .Y(n4498) );
  INVX1 U10953 ( .A(M1_b_14_), .Y(n4502) );
  NAND2X4 U10954 ( .A(n4503), .B(n13261), .Y(n14208) );
  XNOR2X1 U10955 ( .A(n3108), .B(n3204), .Y(n6008) );
  NAND2X1 U10956 ( .A(n18917), .B(n4507), .Y(n18924) );
  NAND3BX2 U10957 ( .AN(n5033), .B(n5472), .C(n4508), .Y(n5888) );
  NAND3X1 U10958 ( .A(n20700), .B(n23734), .C(n4508), .Y(n4887) );
  CLKINVX3 U10959 ( .A(n17493), .Y(n4510) );
  NOR2X1 U10960 ( .A(n4876), .B(n18624), .Y(n6083) );
  XOR2X1 U10961 ( .A(n18603), .B(n3197), .Y(n4876) );
  OAI22X1 U10962 ( .A0(n12635), .A1(n4512), .B0(n12513), .B1(n11670), .Y(
        n11801) );
  XOR2X1 U10963 ( .A(n16884), .B(n4513), .Y(n4512) );
  INVX1 U10964 ( .A(n11791), .Y(n4515) );
  NAND2X4 U10965 ( .A(n4519), .B(n18504), .Y(n18111) );
  NOR2X1 U10966 ( .A(n25813), .B(n2986), .Y(n4521) );
  OAI21X2 U10967 ( .A0(n19014), .A1(n18965), .B0(n18964), .Y(n4523) );
  NOR2X1 U10968 ( .A(n4860), .B(n25900), .Y(n4527) );
  NAND2X1 U10969 ( .A(n25206), .B(data[34]), .Y(n4528) );
  NOR2X1 U10970 ( .A(n15942), .B(n26294), .Y(n4531) );
  NAND2BX4 U10971 ( .AN(n4536), .B(n4535), .Y(M5_b_18_) );
  OAI22X2 U10972 ( .A0(n4541), .A1(n18111), .B0(n18504), .B1(n17621), .Y(
        n17631) );
  OAI22X1 U10973 ( .A0(n4541), .A1(n18504), .B0(n18111), .B1(n17521), .Y(
        n17562) );
  XOR2X1 U10974 ( .A(n3196), .B(n3189), .Y(n4541) );
  NAND2XL U10975 ( .A(n7436), .B(n7435), .Y(n4544) );
  INVX1 U10976 ( .A(n7445), .Y(n7436) );
  NAND3X1 U10977 ( .A(n7442), .B(n7435), .C(n7437), .Y(n4545) );
  AOI21X1 U10978 ( .A0(n25740), .A1(n3065), .B0(n5102), .Y(n5101) );
  NAND2X1 U10979 ( .A(n20882), .B(n3139), .Y(n4546) );
  AOI22X1 U10980 ( .A0(n13463), .A1(n4547), .B0(n13461), .B1(n13462), .Y(
        n13467) );
  AND2X2 U10981 ( .A(n13460), .B(n13459), .Y(n4547) );
  NAND2BX1 U10982 ( .AN(n13461), .B(n4548), .Y(n13463) );
  INVX1 U10983 ( .A(n13462), .Y(n4548) );
  AOI2BB1X2 U10984 ( .A0N(n25731), .A1N(n4582), .B0(n4715), .Y(n4549) );
  NAND3X1 U10985 ( .A(n4551), .B(n11501), .C(n4550), .Y(M1_b_2_) );
  XOR2X2 U10986 ( .A(n4553), .B(n6982), .Y(n6980) );
  NAND2X1 U10987 ( .A(n3139), .B(n23580), .Y(n4555) );
  XNOR2X1 U10988 ( .A(n4556), .B(n9787), .Y(n5745) );
  XNOR2X1 U10989 ( .A(n9788), .B(n4557), .Y(n4556) );
  INVX1 U10990 ( .A(M2_a_14_), .Y(n5761) );
  NAND2X2 U10991 ( .A(n4560), .B(n4559), .Y(n4569) );
  XNOR2X1 U10992 ( .A(M2_a_14_), .B(n10388), .Y(n4560) );
  OAI21X1 U10993 ( .A0(n10656), .A1(n10622), .B0(n10621), .Y(n5227) );
  AOI21X1 U10994 ( .A0(n10627), .A1(n10631), .B0(n10620), .Y(n10621) );
  OAI21X1 U10995 ( .A0(n14585), .A1(n14599), .B0(n14586), .Y(n14000) );
  XNOR2X1 U10996 ( .A(n10324), .B(n10335), .Y(n9272) );
  NAND2X1 U10997 ( .A(n5502), .B(n14533), .Y(n14531) );
  OAI22XL U10998 ( .A0(n18226), .A1(n17866), .B0(n17715), .B1(n18223), .Y(
        n17865) );
  NOR2X1 U10999 ( .A(n5678), .B(n5680), .Y(n5679) );
  OAI21X2 U11000 ( .A0(n13981), .A1(n14400), .B0(n13980), .Y(n5023) );
  XNOR2X1 U11001 ( .A(n14307), .B(n13605), .Y(n13533) );
  NOR2X1 U11002 ( .A(n20929), .B(n3958), .Y(n20346) );
  NOR2X4 U11003 ( .A(n10180), .B(n10186), .Y(n10190) );
  XOR2X1 U11004 ( .A(M2_mult_x_15_n43), .B(n6140), .Y(n6139) );
  OAI22X1 U11005 ( .A0(n11830), .A1(n12222), .B0(n12352), .B1(n6105), .Y(
        n11846) );
  OAI21XL U11006 ( .A0(n25207), .A1(n25206), .B0(n25205), .Y(n25208) );
  AOI22X1 U11007 ( .A0(n24236), .A1(n4215), .B0(n4220), .B1(n24218), .Y(n24226) );
  XNOR2X1 U11008 ( .A(M2_mult_x_15_a_1_), .B(M2_mult_x_15_n1668), .Y(n9301) );
  BUFX3 U11009 ( .A(n9341), .Y(M2_mult_x_15_n1668) );
  NOR2X1 U11010 ( .A(n15150), .B(n15105), .Y(n14786) );
  AOI21XL U11011 ( .A0(n15303), .A1(n3156), .B0(n15313), .Y(n15316) );
  NOR2X1 U11012 ( .A(n5026), .B(n23709), .Y(n5025) );
  OAI21X1 U11013 ( .A0(n6274), .A1(n26218), .B0(n6252), .Y(M0_b_6_) );
  AOI22XL U11014 ( .A0(n6733), .A1(target_temp[6]), .B0(in_valid_d), .B1(w1[6]), .Y(n6252) );
  BUFX3 U11015 ( .A(n5246), .Y(n4811) );
  NAND2X1 U11016 ( .A(n14324), .B(n14323), .Y(n14541) );
  AOI21X1 U11017 ( .A0(n14564), .A1(n14560), .B0(n14522), .Y(n14523) );
  INVX4 U11018 ( .A(n13510), .Y(n14298) );
  NAND2X1 U11019 ( .A(n20282), .B(n20283), .Y(n20365) );
  BUFX4 U11020 ( .A(M0_b_13_), .Y(n25878) );
  BUFX8 U11021 ( .A(n10656), .Y(n5237) );
  AOI21X1 U11022 ( .A0(n10576), .A1(n10562), .B0(n10561), .Y(n10586) );
  AOI22X1 U11023 ( .A0(n4566), .A1(data[20]), .B0(in_valid_d), .B1(w1[276]), 
        .Y(n9063) );
  XNOR2XL U11024 ( .A(M2_a_3_), .B(n10515), .Y(n9383) );
  NOR2BXL U11025 ( .AN(n3110), .B(n16332), .Y(n16608) );
  OAI21XL U11026 ( .A0(n16732), .A1(n16731), .B0(n16730), .Y(n16761) );
  ADDFX2 U11027 ( .A(n25881), .B(n25882), .CI(n7231), .CO(n7303), .S(n7223) );
  XOR2X1 U11028 ( .A(n25881), .B(n26488), .Y(n6487) );
  INVX1 U11029 ( .A(M1_b_6_), .Y(n5152) );
  CLKINVX3 U11030 ( .A(n20810), .Y(n20709) );
  NOR2X2 U11031 ( .A(n10137), .B(n10136), .Y(n10180) );
  OAI22XL U11032 ( .A0(n2997), .A1(n13844), .B0(n13843), .B1(n13842), .Y(
        n13895) );
  NAND2XL U11033 ( .A(n6522), .B(n5553), .Y(n5552) );
  NOR2X1 U11034 ( .A(n6673), .B(n6672), .Y(n6675) );
  XNOR2X1 U11035 ( .A(n7092), .B(n25882), .Y(n6474) );
  NAND2X1 U11036 ( .A(n5770), .B(n4719), .Y(n4825) );
  OAI21XL U11037 ( .A0(n7075), .A1(n7074), .B0(n7073), .Y(n7077) );
  NAND2X1 U11038 ( .A(n5112), .B(n5111), .Y(n6969) );
  AND2X2 U11039 ( .A(n5501), .B(n14543), .Y(n4561) );
  AOI22XL U11040 ( .A0(n25533), .A1(n25664), .B0(n24958), .B1(y11[8]), .Y(
        n24599) );
  XNOR2X1 U11041 ( .A(n9851), .B(n10538), .Y(n9207) );
  CLKINVX3 U11042 ( .A(n14356), .Y(n14353) );
  OR2X2 U11043 ( .A(n6719), .B(n6718), .Y(n6721) );
  ADDFX2 U11044 ( .A(n6430), .B(n6429), .CI(n6428), .CO(n6442), .S(n6466) );
  XNOR2X1 U11045 ( .A(n18500), .B(n3196), .Y(n17746) );
  OAI22X1 U11046 ( .A0(n18226), .A1(n17904), .B0(n17866), .B1(n18223), .Y(
        n17910) );
  NAND3X2 U11047 ( .A(n9071), .B(n5201), .C(n5200), .Y(M2_a_19_) );
  NAND2X2 U11048 ( .A(n9215), .B(n5199), .Y(n10532) );
  CLKINVX3 U11049 ( .A(n6289), .Y(n6744) );
  OAI22XL U11050 ( .A0(n13315), .A1(n13790), .B0(n13390), .B1(n13721), .Y(
        n13376) );
  XNOR2X2 U11051 ( .A(n14628), .B(n14627), .Y(n20982) );
  OAI21XL U11052 ( .A0(n14638), .A1(n14624), .B0(n14623), .Y(n14628) );
  NAND2X1 U11053 ( .A(n5100), .B(n20894), .Y(n20895) );
  OAI21X1 U11054 ( .A0(n6274), .A1(n26215), .B0(n6248), .Y(M0_b_11_) );
  OAI21X2 U11055 ( .A0(n7382), .A1(n26011), .B0(n2994), .Y(n6288) );
  XNOR2X1 U11056 ( .A(M5_mult_x_15_n1), .B(n3196), .Y(n16335) );
  AOI21X1 U11057 ( .A0(n14496), .A1(n14495), .B0(n14494), .Y(n14497) );
  NAND2X1 U11058 ( .A(n14689), .B(n14688), .Y(n14690) );
  OAI21X2 U11059 ( .A0(n7382), .A1(n25999), .B0(n6247), .Y(M0_a_7_) );
  AOI21X4 U11060 ( .A0(n7672), .A1(n7782), .B0(n7671), .Y(n7822) );
  INVX1 U11061 ( .A(n7782), .Y(n7757) );
  OAI21X2 U11062 ( .A0(n7490), .A1(n7489), .B0(n7488), .Y(n7782) );
  INVX1 U11063 ( .A(n6298), .Y(n7556) );
  AOI21X1 U11064 ( .A0(n4635), .A1(n6664), .B0(n6663), .Y(n5555) );
  AND2X2 U11065 ( .A(n6660), .B(n6659), .Y(n6664) );
  OAI22XL U11066 ( .A0(n6845), .A1(n6605), .B0(n6604), .B1(n6843), .Y(n6611)
         );
  XNOR2X1 U11067 ( .A(n21054), .B(n7475), .Y(n6516) );
  XNOR2X1 U11068 ( .A(n21054), .B(M0_b_11_), .Y(n6471) );
  INVX1 U11069 ( .A(n6231), .Y(n25871) );
  ADDFX2 U11070 ( .A(n6940), .B(n6939), .CI(n6938), .CO(n6984), .S(n6936) );
  ADDFX2 U11071 ( .A(n18607), .B(n18606), .CI(n18605), .CO(n18627), .S(n18613)
         );
  OAI22X1 U11072 ( .A0(n18659), .A1(n18482), .B0(n17832), .B1(n18609), .Y(
        n18606) );
  NAND2X1 U11073 ( .A(n4579), .B(w1[18]), .Y(n5132) );
  OAI22X1 U11074 ( .A0(n17148), .A1(M3_mult_x_15_b_9_), .B0(n3194), .B1(n16884), .Y(n6013) );
  ADDFX2 U11075 ( .A(n16884), .B(n3190), .CI(n16872), .CO(n16886), .S(n16934)
         );
  NOR2X2 U11076 ( .A(n5917), .B(n3121), .Y(n25638) );
  INVX4 U11077 ( .A(n5374), .Y(n18428) );
  ADDFX2 U11078 ( .A(n10025), .B(n10024), .CI(n10023), .CO(n10015), .S(n10026)
         );
  OAI22XL U11079 ( .A0(n9966), .A1(n9964), .B0(n10159), .B1(n9817), .Y(n9955)
         );
  OAI22X1 U11080 ( .A0(n4642), .A1(n7297), .B0(n7465), .B1(n7712), .Y(n7474)
         );
  OAI21X1 U11081 ( .A0(n7670), .A1(n7754), .B0(n7669), .Y(n7671) );
  NOR2X2 U11082 ( .A(n7670), .B(n7752), .Y(n7672) );
  OAI22X1 U11083 ( .A0(n7292), .A1(n5124), .B0(n7695), .B1(n7467), .Y(n7463)
         );
  XOR2X2 U11084 ( .A(n18833), .B(n18794), .Y(n24250) );
  OAI22XL U11085 ( .A0(n18083), .A1(n18000), .B0(n18429), .B1(n17974), .Y(
        n18018) );
  OAI22X1 U11086 ( .A0(n17092), .A1(n6014), .B0(n16317), .B1(n16013), .Y(
        n16070) );
  OAI21X1 U11087 ( .A0(n25731), .A1(n3024), .B0(n25005), .Y(n5001) );
  OAI22X1 U11088 ( .A0(n10517), .A1(n9398), .B0(n10533), .B1(n9318), .Y(n9425)
         );
  OAI21X1 U11089 ( .A0(n3494), .A1(n7748), .B0(n7747), .Y(n7751) );
  NOR2X1 U11090 ( .A(n23743), .B(n5387), .Y(n5386) );
  NAND2BX1 U11091 ( .AN(n20667), .B(n23744), .Y(n5026) );
  NOR2X4 U11092 ( .A(in_valid_t), .B(n25693), .Y(n11481) );
  NAND2X1 U11093 ( .A(n12510), .B(n12509), .Y(n12915) );
  INVX4 U11094 ( .A(n21166), .Y(n15941) );
  OAI22X1 U11095 ( .A0(n12717), .A1(n11762), .B0(n12718), .B1(n11877), .Y(
        n11883) );
  XNOR2X1 U11096 ( .A(n12716), .B(n3190), .Y(n11762) );
  ADDFX2 U11097 ( .A(n13683), .B(n13682), .CI(n13681), .CO(n13739), .S(n13749)
         );
  NOR2X1 U11098 ( .A(n4821), .B(n4819), .Y(n23547) );
  AOI22X2 U11099 ( .A0(n23539), .A1(n3455), .B0(n23611), .B1(n3139), .Y(n23604) );
  XOR2X1 U11100 ( .A(n20818), .B(n20817), .Y(n23539) );
  OAI22X1 U11101 ( .A0(n7287), .A1(n6929), .B0(n6976), .B1(n7288), .Y(n6975)
         );
  AOI22X2 U11102 ( .A0(n20939), .A1(n5336), .B0(n20938), .B1(n3136), .Y(n24249) );
  OAI21X1 U11103 ( .A0(n3494), .A1(n7685), .B0(n7684), .Y(n7700) );
  XNOR2X1 U11104 ( .A(n3209), .B(n7569), .Y(n6365) );
  NAND2X1 U11105 ( .A(n9089), .B(n11533), .Y(M2_b_16_) );
  XNOR2X1 U11106 ( .A(n9851), .B(n10335), .Y(n9320) );
  AOI21X1 U11107 ( .A0(n14606), .A1(n14626), .B0(n14605), .Y(n14607) );
  OAI22X1 U11108 ( .A0(n13790), .A1(n25860), .B0(n13721), .B1(n13720), .Y(
        n13775) );
  OAI22X1 U11109 ( .A0(n9504), .A1(n9460), .B0(n10496), .B1(n9505), .Y(n9514)
         );
  NAND2X1 U11110 ( .A(n10143), .B(n10142), .Y(n10238) );
  NOR2X1 U11111 ( .A(n18688), .B(n18687), .Y(n18951) );
  AOI21X1 U11112 ( .A0(n18690), .A1(n18934), .B0(n18689), .Y(n18691) );
  ADDFX2 U11113 ( .A(n7161), .B(n7160), .CI(n7159), .CO(n7178), .S(n7140) );
  AOI222X1 U11114 ( .A0(n23721), .A1(n25737), .B0(n25743), .B1(y20[17]), .C0(
        n25422), .C1(n20890), .Y(n2377) );
  NAND2X1 U11115 ( .A(n10067), .B(n10065), .Y(n4562) );
  NAND2X1 U11116 ( .A(n10066), .B(n10065), .Y(n4563) );
  NAND3X1 U11117 ( .A(n4564), .B(n4562), .C(n4563), .Y(n10059) );
  XNOR2X1 U11118 ( .A(n5745), .B(n5177), .Y(n5176) );
  NOR2X4 U11119 ( .A(n10213), .B(n10208), .Y(n10135) );
  AOI22XL U11120 ( .A0(n11536), .A1(data[1]), .B0(in_valid_d), .B1(w1[257]), 
        .Y(n9096) );
  NAND2X2 U11121 ( .A(n14550), .B(n14322), .Y(n14532) );
  XNOR2X1 U11122 ( .A(M2_mult_x_15_a_1_), .B(n10386), .Y(n9736) );
  NOR2X2 U11123 ( .A(n10476), .B(n10475), .Y(n10623) );
  NOR2BX2 U11124 ( .AN(n10580), .B(n5007), .Y(n5006) );
  OAI22X1 U11125 ( .A0(n10517), .A1(n10366), .B0(n10533), .B1(n10380), .Y(
        n10391) );
  XNOR2X1 U11126 ( .A(n10494), .B(n10538), .Y(n10380) );
  NAND2X4 U11127 ( .A(n9203), .B(n10369), .Y(n10368) );
  XNOR2X2 U11128 ( .A(n14635), .B(n14634), .Y(n23589) );
  BUFX3 U11129 ( .A(M1_a_7_), .Y(n14027) );
  INVX1 U11130 ( .A(n24984), .Y(n25753) );
  INVXL U11131 ( .A(n14080), .Y(n6056) );
  OAI21XL U11132 ( .A0(n24656), .A1(n3121), .B0(n23913), .Y(n2594) );
  XOR2X1 U11133 ( .A(n23649), .B(n23648), .Y(n23792) );
  ADDFX2 U11134 ( .A(n9535), .B(n9534), .CI(n9533), .CO(n9569), .S(n9553) );
  XNOR2X2 U11135 ( .A(n14518), .B(n14517), .Y(n14683) );
  XOR2X2 U11136 ( .A(n5092), .B(n14642), .Y(n23588) );
  XNOR2X1 U11137 ( .A(n10339), .B(n10311), .Y(n9382) );
  XNOR2X2 U11138 ( .A(n14531), .B(n14530), .Y(n14685) );
  OAI22XL U11139 ( .A0(n9983), .A1(n9815), .B0(n9981), .B1(n9785), .Y(n9821)
         );
  XNOR2X1 U11140 ( .A(n9904), .B(n10342), .Y(n9785) );
  XNOR2X1 U11141 ( .A(n25885), .B(n9863), .Y(n9266) );
  NOR2X2 U11142 ( .A(n5275), .B(n20972), .Y(n5274) );
  OAI22X1 U11143 ( .A0(n10368), .A1(n9265), .B0(n10369), .B1(n9264), .Y(n9277)
         );
  XNOR2X2 U11144 ( .A(n14566), .B(n14565), .Y(n14687) );
  OAI22XL U11145 ( .A0(n13556), .A1(n13721), .B0(n13538), .B1(n13790), .Y(
        n13574) );
  OAI22X1 U11146 ( .A0(n13650), .A1(n13721), .B0(n13620), .B1(n13790), .Y(
        n13659) );
  OAI22XL U11147 ( .A0(n13860), .A1(n14044), .B0(n13872), .B1(n13974), .Y(
        n13894) );
  AND4X4 U11148 ( .A(n14684), .B(n23745), .C(n14682), .D(n14683), .Y(n6072) );
  OAI22XL U11149 ( .A0(n9966), .A1(n9753), .B0(n10159), .B1(n9728), .Y(n9758)
         );
  OAI22X1 U11150 ( .A0(n9445), .A1(n9614), .B0(n9906), .B1(n9444), .Y(n9605)
         );
  OAI22X1 U11151 ( .A0(n13367), .A1(n14198), .B0(n13363), .B1(n14208), .Y(
        n13365) );
  XNOR2X1 U11152 ( .A(n13864), .B(M1_b_15_), .Y(n13363) );
  OAI22XL U11153 ( .A0(n13652), .A1(n2997), .B0(n13701), .B1(n13843), .Y(
        n13675) );
  OAI22XL U11154 ( .A0(n9551), .A1(n9771), .B0(n9974), .B1(n9735), .Y(n9776)
         );
  OAI22X1 U11155 ( .A0(n10368), .A1(n9773), .B0(n9780), .B1(n9772), .Y(n9794)
         );
  OAI22X1 U11156 ( .A0(n9963), .A1(n9631), .B0(n9595), .B1(n3180), .Y(n9634)
         );
  XNOR2XL U11157 ( .A(n25864), .B(n23173), .Y(n14209) );
  AOI21X1 U11158 ( .A0(n14427), .A1(y10[6]), .B0(n5346), .Y(n5345) );
  XNOR2X1 U11159 ( .A(M2_mult_x_15_a_1_), .B(M2_b_15_), .Y(n9693) );
  XNOR2X1 U11160 ( .A(M2_mult_x_15_n43), .B(M2_b_15_), .Y(n9502) );
  XNOR2X1 U11161 ( .A(n9851), .B(M2_b_15_), .Y(n9421) );
  XNOR2X1 U11162 ( .A(n10324), .B(M2_b_15_), .Y(n9226) );
  XNOR2X1 U11163 ( .A(n9904), .B(M2_b_15_), .Y(n9640) );
  NAND2X4 U11164 ( .A(n9088), .B(n11527), .Y(M2_b_15_) );
  OAI22X1 U11165 ( .A0(n13284), .A1(n14080), .B0(n13283), .B1(n3173), .Y(
        n13288) );
  OAI22XL U11166 ( .A0(n13328), .A1(n13606), .B0(n13391), .B1(n3181), .Y(
        n13373) );
  XNOR2X1 U11167 ( .A(n14195), .B(n13693), .Y(n13315) );
  OAI22X1 U11168 ( .A0(n13266), .A1(n14029), .B0(n13219), .B1(n14044), .Y(
        n13291) );
  OAI22XL U11169 ( .A0(n9979), .A1(n9755), .B0(n9977), .B1(n9734), .Y(n9777)
         );
  OAI22XL U11170 ( .A0(n14080), .A1(n25861), .B0(n3173), .B1(n5489), .Y(n14090) );
  XNOR2X1 U11171 ( .A(n14236), .B(n14228), .Y(n13963) );
  XNOR2X1 U11172 ( .A(n14236), .B(n4848), .Y(n13446) );
  XNOR2XL U11173 ( .A(n14236), .B(n13204), .Y(n13282) );
  OAI22XL U11174 ( .A0(n9963), .A1(n9301), .B0(n3180), .B1(M2_mult_x_15_a_1_), 
        .Y(n9305) );
  OAI21X1 U11175 ( .A0(n6274), .A1(n26228), .B0(n6237), .Y(M0_b_17_) );
  OAI22XL U11176 ( .A0(n13286), .A1(n13721), .B0(n13218), .B1(n13790), .Y(
        n13292) );
  OAI22X1 U11177 ( .A0(n9966), .A1(n9728), .B0(n10159), .B1(n9699), .Y(n9733)
         );
  OAI211X2 U11178 ( .A0(n25915), .A1(n3103), .B0(n9094), .C0(n9093), .Y(
        M2_a_22_) );
  AND2X2 U11179 ( .A(n4566), .B(learning_rate[13]), .Y(n5513) );
  XNOR2X1 U11180 ( .A(n9851), .B(n10539), .Y(n9227) );
  AOI22X1 U11181 ( .A0(n4566), .A1(data[15]), .B0(in_valid_d), .B1(w1[271]), 
        .Y(n9088) );
  OAI22XL U11182 ( .A0(n9963), .A1(n9782), .B0(n9736), .B1(n3180), .Y(n9779)
         );
  INVX8 U11183 ( .A(n13280), .Y(n14198) );
  OAI22X1 U11184 ( .A0(n13914), .A1(n14208), .B0(n13976), .B1(n14198), .Y(
        n13961) );
  OAI22X1 U11185 ( .A0(n10296), .A1(n9774), .B0(n9959), .B1(n9729), .Y(n9757)
         );
  OAI21XL U11186 ( .A0(n24697), .A1(n3121), .B0(n23902), .Y(n2590) );
  NAND2X1 U11187 ( .A(n9073), .B(n11511), .Y(M2_b_6_) );
  OAI22X1 U11188 ( .A0(n13653), .A1(n14208), .B0(n13700), .B1(n14198), .Y(
        n13674) );
  INVX4 U11189 ( .A(n13258), .Y(n14157) );
  NOR2X1 U11190 ( .A(n25755), .B(n25255), .Y(n25760) );
  OAI22X1 U11191 ( .A0(n13861), .A1(n14157), .B0(n13876), .B1(n14120), .Y(
        n13893) );
  XNOR2X1 U11192 ( .A(n9851), .B(n9839), .Y(n9771) );
  INVX8 U11193 ( .A(in_valid_d), .Y(n4581) );
  INVX8 U11194 ( .A(in_valid_d), .Y(n4582) );
  INVX8 U11195 ( .A(in_valid_d), .Y(n4583) );
  INVX8 U11196 ( .A(in_valid_d), .Y(n4584) );
  INVX8 U11197 ( .A(in_valid_d), .Y(n4586) );
  INVXL U11198 ( .A(n8524), .Y(n8339) );
  CLKINVX3 U11199 ( .A(n21055), .Y(n10295) );
  INVXL U11200 ( .A(n4565), .Y(n14062) );
  OAI22XL U11201 ( .A0(n14044), .A1(n14030), .B0(n14029), .B1(n6210), .Y(
        n14060) );
  NAND2X1 U11202 ( .A(n6152), .B(n5240), .Y(n5239) );
  XOR2XL U11203 ( .A(M2_a_18_), .B(M2_a_19_), .Y(n5199) );
  OAI21XL U11204 ( .A0(n15013), .A1(n15012), .B0(n15011), .Y(n15014) );
  OAI21X1 U11205 ( .A0(n17167), .A1(n26003), .B0(n4894), .Y(n5971) );
  NAND2X1 U11206 ( .A(n4826), .B(target_temp[20]), .Y(n11543) );
  NOR2XL U11207 ( .A(n11691), .B(n12338), .Y(n11645) );
  OAI22XL U11208 ( .A0(n12995), .A1(M3_mult_x_15_b_3_), .B0(n12535), .B1(
        n12271), .Y(n11657) );
  AOI21XL U11209 ( .A0(n23001), .A1(n11071), .B0(n22969), .Y(n22655) );
  AND2X2 U11210 ( .A(in_valid_t), .B(w2[11]), .Y(n4655) );
  OAI22X1 U11211 ( .A0(n5455), .A1(n17832), .B0(n17637), .B1(n18659), .Y(
        n17732) );
  OAI22XL U11212 ( .A0(n18652), .A1(n17638), .B0(n17872), .B1(n17745), .Y(
        n17731) );
  OAI2BB1XL U11213 ( .A0N(n6123), .A1N(n17624), .B0(n6122), .Y(n17736) );
  OAI22XL U11214 ( .A0(n5893), .A1(n17750), .B0(n17623), .B1(n18541), .Y(
        n17737) );
  OAI21XL U11215 ( .A0(n7822), .A1(n7683), .B0(n7682), .Y(n7704) );
  NAND4XL U11216 ( .A(n20161), .B(n24716), .C(n24680), .D(n24798), .Y(n20162)
         );
  NOR2XL U11217 ( .A(n20160), .B(n20159), .Y(n20161) );
  NAND4XL U11218 ( .A(n20158), .B(n20236), .C(n20195), .D(n20196), .Y(n20159)
         );
  NAND3XL U11219 ( .A(n20235), .B(n20186), .C(n20188), .Y(n20160) );
  NAND2XL U11220 ( .A(n19978), .B(n19977), .Y(n19979) );
  INVXL U11221 ( .A(n19976), .Y(n19978) );
  NAND2XL U11222 ( .A(n19973), .B(n19972), .Y(n19974) );
  INVXL U11223 ( .A(n19971), .Y(n19973) );
  NAND2XL U11224 ( .A(n20007), .B(n20005), .Y(n19969) );
  INVXL U11225 ( .A(n20004), .Y(n19967) );
  AND4XL U11226 ( .A(n24275), .B(n20795), .C(n24348), .D(n20787), .Y(n18969)
         );
  NAND2XL U11227 ( .A(n22165), .B(n22167), .Y(n22139) );
  INVXL U11228 ( .A(n22138), .Y(n22140) );
  AOI31XL U11229 ( .A0(n22156), .A1(n22137), .A2(n22160), .B0(n22136), .Y(
        n22138) );
  NAND3BXL U11230 ( .AN(n7874), .B(n23850), .C(n23683), .Y(n7875) );
  INVXL U11231 ( .A(n23685), .Y(n7876) );
  NAND4XL U11232 ( .A(n23854), .B(n23822), .C(n23865), .D(n23782), .Y(n7874)
         );
  NAND4XL U11233 ( .A(n14426), .B(n14425), .C(n14424), .D(n14423), .Y(n14428)
         );
  NAND4XL U11234 ( .A(n14422), .B(n14421), .C(n14420), .D(n14419), .Y(n14429)
         );
  NOR4XL U11235 ( .A(n20795), .B(n24348), .C(n20787), .D(n20786), .Y(n18789)
         );
  INVXL U11236 ( .A(n24275), .Y(n18787) );
  NAND2XL U11237 ( .A(n8977), .B(n8979), .Y(n8951) );
  INVXL U11238 ( .A(n8950), .Y(n8952) );
  AOI31XL U11239 ( .A0(n8968), .A1(n8949), .A2(n8972), .B0(n8948), .Y(n8950)
         );
  XOR2XL U11240 ( .A(n22705), .B(n3058), .Y(n23048) );
  NAND2XL U11241 ( .A(n22928), .B(n22987), .Y(n4706) );
  NAND2BXL U11242 ( .AN(n6944), .B(n4789), .Y(n6480) );
  AOI22X1 U11243 ( .A0(n4566), .A1(data[11]), .B0(in_valid_d), .B1(w1[267]), 
        .Y(n9049) );
  XNOR2XL U11244 ( .A(n14235), .B(n25861), .Y(n13714) );
  AOI2BB2XL U11245 ( .B0(n8514), .B1(n3087), .A0N(n8434), .A1N(n8431), .Y(
        n8432) );
  OAI21XL U11246 ( .A0(n3162), .A1(n8380), .B0(n8344), .Y(n8406) );
  AOI222XL U11247 ( .A0(n22988), .A1(n10769), .B0(n22980), .B1(n23002), .C0(
        n22976), .C1(n10749), .Y(n22915) );
  CMPR32X1 U11248 ( .A(n6530), .B(n6529), .C(n6528), .CO(n6677), .S(n6688) );
  OAI21XL U11249 ( .A0(n6274), .A1(n26225), .B0(n6270), .Y(n6830) );
  AOI22X1 U11250 ( .A0(n7389), .A1(target_temp[16]), .B0(n3123), .B1(w1[16]), 
        .Y(n6270) );
  INVX8 U11251 ( .A(n10295), .Y(n10324) );
  CLKINVX2 U11252 ( .A(M2_a_17_), .Y(n5202) );
  AOI22X1 U11253 ( .A0(n9164), .A1(y12[7]), .B0(n14427), .B1(y10[7]), .Y(n9066) );
  NAND2X1 U11254 ( .A(n4856), .B(y12[6]), .Y(n5344) );
  NOR2X1 U11255 ( .A(n3103), .B(n25912), .Y(n5080) );
  INVXL U11256 ( .A(M2_mult_x_15_a_1_), .Y(n9222) );
  CLKINVX3 U11257 ( .A(n5489), .Y(n25861) );
  NOR2XL U11258 ( .A(n25860), .B(n23174), .Y(M1_U4_U1_or2_tree_0__1__28_) );
  NAND2X1 U11259 ( .A(in_valid_d), .B(w1[140]), .Y(n5342) );
  NAND2X1 U11260 ( .A(in_valid_d), .B(w1[141]), .Y(n6086) );
  OAI21XL U11261 ( .A0(n25243), .A1(n25912), .B0(n9042), .Y(M1_a_20_) );
  BUFX3 U11262 ( .A(M1_a_19_), .Y(n14288) );
  INVX1 U11263 ( .A(n23123), .Y(n21445) );
  OAI21XL U11264 ( .A0(n14967), .A1(n15074), .B0(n15073), .Y(n15394) );
  OAI211XL U11265 ( .A0(n3090), .A1(n15236), .B0(n15046), .C0(n15072), .Y(
        n15074) );
  NAND2XL U11266 ( .A(n15224), .B(n3090), .Y(n15072) );
  INVXL U11267 ( .A(n22947), .Y(n22959) );
  AOI222XL U11268 ( .A0(n23152), .A1(n23002), .B0(n23093), .B1(n10749), .C0(
        n23150), .C1(n3116), .Y(n22946) );
  XOR2XL U11269 ( .A(n22922), .B(n3056), .Y(M6_mult_x_15_n1102) );
  XOR2XL U11270 ( .A(n22934), .B(n3053), .Y(M6_mult_x_15_n1174) );
  XOR2XL U11271 ( .A(n21090), .B(n21089), .Y(M6_mult_x_15_n1126) );
  XOR2XL U11272 ( .A(n22721), .B(n3058), .Y(n23031) );
  AOI222XL U11273 ( .A0(n22928), .A1(n10769), .B0(n22700), .B1(n23002), .C0(
        n22927), .C1(n10749), .Y(n22720) );
  XOR2XL U11274 ( .A(n22648), .B(n22647), .Y(n23142) );
  NAND2XL U11275 ( .A(n22646), .B(n22645), .Y(n22647) );
  INVXL U11276 ( .A(n22644), .Y(n22646) );
  XOR2XL U11277 ( .A(n22707), .B(n3119), .Y(n23047) );
  AOI222XL U11278 ( .A0(n22892), .A1(n10749), .B0(n22708), .B1(n3116), .C0(
        n22891), .C1(n22987), .Y(n22706) );
  CLKINVX3 U11279 ( .A(n26495), .Y(n26496) );
  INVXL U11280 ( .A(n11165), .Y(n10770) );
  AOI21XL U11281 ( .A0(n22952), .A1(n11071), .B0(n10797), .Y(n22681) );
  NOR2X1 U11282 ( .A(n17167), .B(n25922), .Y(n5680) );
  NOR2X1 U11283 ( .A(n4860), .B(n26020), .Y(n5678) );
  NAND2XL U11284 ( .A(n21166), .B(target_temp[3]), .Y(n4753) );
  AOI22X1 U11285 ( .A0(n25229), .A1(y12[22]), .B0(n14427), .B1(y10[22]), .Y(
        n9094) );
  OAI22X1 U11286 ( .A0(n12618), .A1(n11816), .B0(n12119), .B1(n11743), .Y(
        n11835) );
  XNOR2XL U11287 ( .A(n12233), .B(n3021), .Y(n11746) );
  BUFX3 U11288 ( .A(M3_mult_x_15_b_13_), .Y(n12560) );
  INVXL U11289 ( .A(M1_b_22_), .Y(n13609) );
  BUFX3 U11290 ( .A(n16319), .Y(n16375) );
  NOR2XL U11291 ( .A(M4_U3_U1_or2_inv_0__30_), .B(n18223), .Y(n17514) );
  OAI21X1 U11292 ( .A0(n17512), .A1(n12271), .B0(n5028), .Y(n17515) );
  AOI21XL U11293 ( .A0(n8673), .A1(n8823), .B0(n3155), .Y(n8672) );
  OAI211XL U11294 ( .A0(n3154), .A1(n8671), .B0(n8295), .C0(n8670), .Y(n8673)
         );
  AOI21XL U11295 ( .A0(n19507), .A1(n19952), .B0(n3164), .Y(n19506) );
  OAI21XL U11296 ( .A0(n3165), .A1(n19550), .B0(n19549), .Y(n19765) );
  AOI21XL U11297 ( .A0(n19550), .A1(n19952), .B0(n3164), .Y(n19549) );
  OAI211XL U11298 ( .A0(n3090), .A1(n15252), .B0(n15046), .C0(n15094), .Y(
        n15096) );
  NAND2XL U11299 ( .A(n15244), .B(n3090), .Y(n15094) );
  NOR2X1 U11300 ( .A(n23402), .B(n21445), .Y(n21478) );
  NAND2XL U11301 ( .A(n21329), .B(temp0[7]), .Y(n21211) );
  NAND2XL U11302 ( .A(n21331), .B(temp0[12]), .Y(n21236) );
  NAND2XL U11303 ( .A(n21331), .B(temp0[11]), .Y(n21238) );
  OAI21XL U11304 ( .A0(n14967), .A1(n15125), .B0(n15124), .Y(n15386) );
  AOI22XL U11305 ( .A0(n15122), .A1(n15121), .B0(n15355), .B1(n15554), .Y(
        n15123) );
  OAI21XL U11306 ( .A0(n14967), .A1(n15168), .B0(n15167), .Y(n15384) );
  NAND2XL U11307 ( .A(n15166), .B(n15256), .Y(n15168) );
  AOI22XL U11308 ( .A0(n15165), .A1(n15355), .B0(n15164), .B1(n15340), .Y(
        n15166) );
  XOR2X2 U11309 ( .A(n3200), .B(n17038), .Y(n16319) );
  ADDFX2 U11310 ( .A(n5430), .B(M3_mult_x_15_b_9_), .CI(n16963), .CO(n16985), 
        .S(n16989) );
  XNOR2XL U11311 ( .A(n22559), .B(n22558), .Y(n23101) );
  NAND2XL U11312 ( .A(n22557), .B(n22556), .Y(n22558) );
  AOI21XL U11313 ( .A0(n22570), .A1(n22568), .B0(n22554), .Y(n22559) );
  INVXL U11314 ( .A(n22555), .Y(n22557) );
  OAI22XL U11315 ( .A0(n17551), .A1(n18541), .B0(n5893), .B1(n17510), .Y(
        n17499) );
  INVX4 U11316 ( .A(n18637), .Y(n18638) );
  XOR3X2 U11317 ( .A(n16394), .B(n16395), .C(n16393), .Y(n16455) );
  NOR2X1 U11318 ( .A(n15940), .B(n25931), .Y(n5648) );
  NOR2X1 U11319 ( .A(n15942), .B(n26296), .Y(n5649) );
  OAI22X1 U11320 ( .A0(n6205), .A1(n15942), .B0(n25914), .B1(n25796), .Y(
        n11487) );
  NAND2X1 U11321 ( .A(in_valid_t), .B(learning_rate[10]), .Y(n6148) );
  NAND2X2 U11322 ( .A(n11628), .B(n5416), .Y(n12578) );
  NAND2XL U11323 ( .A(n8698), .B(n8697), .Y(n8745) );
  INVXL U11324 ( .A(n8781), .Y(n8860) );
  NAND2XL U11325 ( .A(n15445), .B(n15444), .Y(n15499) );
  INVXL U11326 ( .A(n22093), .Y(n22128) );
  NAND2XL U11327 ( .A(n21329), .B(temp0[8]), .Y(n21209) );
  NOR2XL U11328 ( .A(n4623), .B(n22186), .Y(n22131) );
  XOR2XL U11329 ( .A(n22120), .B(n22119), .Y(n22295) );
  NAND2XL U11330 ( .A(n6202), .B(n22118), .Y(n22119) );
  XOR2XL U11331 ( .A(n22110), .B(n22109), .Y(n22292) );
  NAND2XL U11332 ( .A(n22108), .B(n22107), .Y(n22109) );
  INVXL U11333 ( .A(n22106), .Y(n22108) );
  NAND2X1 U11334 ( .A(n4875), .B(n4721), .Y(n5411) );
  NAND2XL U11335 ( .A(n11108), .B(n10938), .Y(n10940) );
  AOI21XL U11336 ( .A0(n11107), .A1(n10938), .B0(n10937), .Y(n10939) );
  NOR2XL U11337 ( .A(n11119), .B(n11109), .Y(n10938) );
  INVXL U11338 ( .A(n7822), .Y(n7793) );
  NAND2XL U11339 ( .A(n19894), .B(n19893), .Y(n19895) );
  INVXL U11340 ( .A(n19892), .Y(n19894) );
  NAND2XL U11341 ( .A(n15495), .B(n15494), .Y(n15496) );
  INVXL U11342 ( .A(n15490), .Y(n15493) );
  NAND2XL U11343 ( .A(n15487), .B(n15486), .Y(n15488) );
  INVXL U11344 ( .A(n15485), .Y(n15487) );
  NAND2XL U11345 ( .A(n15594), .B(n15593), .Y(n15595) );
  INVXL U11346 ( .A(n15592), .Y(n15594) );
  NAND2XL U11347 ( .A(n15616), .B(n15615), .Y(n15617) );
  INVXL U11348 ( .A(n15614), .Y(n15616) );
  NAND2XL U11349 ( .A(n21954), .B(n21953), .Y(n21955) );
  AOI21XL U11350 ( .A0(n22117), .A1(n21951), .B0(n21950), .Y(n21956) );
  INVXL U11351 ( .A(n21952), .Y(n21954) );
  NAND2XL U11352 ( .A(n21945), .B(n21944), .Y(n21946) );
  INVXL U11353 ( .A(n21943), .Y(n21945) );
  NAND2XL U11354 ( .A(n21940), .B(n21939), .Y(n21941) );
  INVXL U11355 ( .A(n21938), .Y(n21940) );
  NAND2XL U11356 ( .A(n15628), .B(n15626), .Y(n15590) );
  INVXL U11357 ( .A(n15625), .Y(n15588) );
  NAND2XL U11358 ( .A(n15622), .B(n15621), .Y(n15623) );
  NAND2BXL U11359 ( .AN(n20637), .B(n9195), .Y(n10287) );
  NOR3XL U11360 ( .A(n23662), .B(n23661), .C(n9194), .Y(n9195) );
  NAND3BXL U11361 ( .AN(n24383), .B(n9193), .C(n24267), .Y(n9194) );
  NOR2XL U11362 ( .A(n25775), .B(n14472), .Y(n14473) );
  NOR4XL U11363 ( .A(n24410), .B(n24083), .C(n24331), .D(n24304), .Y(n14471)
         );
  INVXL U11364 ( .A(n24280), .Y(n14469) );
  NAND3BXL U11365 ( .AN(n14655), .B(n25774), .C(n24105), .Y(n14656) );
  INVXL U11366 ( .A(n25775), .Y(n14657) );
  NAND4XL U11367 ( .A(n24280), .B(n24410), .C(n24083), .D(n24331), .Y(n14655)
         );
  INVXL U11368 ( .A(n20115), .Y(n20116) );
  NAND2XL U11369 ( .A(n20114), .B(n20113), .Y(n20118) );
  NAND2XL U11370 ( .A(n3126), .B(n22305), .Y(n22235) );
  OAI21XL U11371 ( .A0(n21365), .A1(n21364), .B0(n21363), .Y(n21389) );
  AOI21XL U11372 ( .A0(n21349), .A1(n21348), .B0(n21347), .Y(n21365) );
  OAI22XL U11373 ( .A0(n22426), .A1(n22317), .B0(n22316), .B1(n3129), .Y(
        n22361) );
  NAND2XL U11374 ( .A(n3126), .B(n22421), .Y(n22257) );
  NOR2XL U11375 ( .A(n22425), .B(n22424), .Y(n22454) );
  NOR2XL U11376 ( .A(n22308), .B(n22423), .Y(n22424) );
  NOR2XL U11377 ( .A(n3126), .B(n22422), .Y(n22425) );
  INVXL U11378 ( .A(n22421), .Y(n22422) );
  INVXL U11379 ( .A(n22165), .Y(n22166) );
  NAND2XL U11380 ( .A(n22164), .B(n22163), .Y(n22168) );
  OAI31XL U11381 ( .A0(n22282), .A1(n22285), .A2(n22162), .B0(n22161), .Y(
        n22163) );
  NAND2XL U11382 ( .A(n4826), .B(target_temp[24]), .Y(n14452) );
  NOR4XL U11383 ( .A(n25181), .B(n25099), .C(n24360), .D(n24359), .Y(n17199)
         );
  INVXL U11384 ( .A(n25107), .Y(n17197) );
  XOR2XL U11385 ( .A(n9149), .B(n10678), .Y(n9169) );
  NAND2XL U11386 ( .A(n20576), .B(n20517), .Y(n20590) );
  OAI21XL U11387 ( .A0(n26282), .A1(n3115), .B0(n14408), .Y(n14698) );
  AOI21XL U11388 ( .A0(y11[24]), .A1(n14417), .B0(n25218), .Y(n14408) );
  XOR2XL U11389 ( .A(n18764), .B(n19035), .Y(n18775) );
  NOR2X1 U11390 ( .A(n3143), .B(n24026), .Y(n4842) );
  NAND2BXL U11391 ( .AN(n24025), .B(n24029), .Y(n24026) );
  NOR2BXL U11392 ( .AN(n20129), .B(n24301), .Y(n20132) );
  OAI22XL U11393 ( .A0(n22267), .A1(n22124), .B0(n22239), .B1(n3082), .Y(
        n22380) );
  NAND2X1 U11394 ( .A(n22359), .B(n3079), .Y(n22389) );
  NAND2XL U11395 ( .A(n23242), .B(n23265), .Y(n22391) );
  NAND2XL U11396 ( .A(n3082), .B(n22392), .Y(n22462) );
  AND4XL U11397 ( .A(n25107), .B(n25181), .C(n25099), .D(n24360), .Y(n17201)
         );
  NAND2XL U11398 ( .A(n3123), .B(w1[151]), .Y(n14453) );
  NAND2XL U11399 ( .A(n25233), .B(learning_rate[23]), .Y(n14454) );
  NAND4XL U11400 ( .A(n14456), .B(n14452), .C(n14451), .D(n14450), .Y(n14714)
         );
  NAND2XL U11401 ( .A(in_valid_d), .B(w1[152]), .Y(n14450) );
  NAND2XL U11402 ( .A(n25233), .B(learning_rate[24]), .Y(n14451) );
  NAND2XL U11403 ( .A(in_valid_d), .B(w1[154]), .Y(n14442) );
  NAND2XL U11404 ( .A(n25233), .B(learning_rate[26]), .Y(n14443) );
  NOR2XL U11405 ( .A(n18786), .B(n18783), .Y(n13021) );
  NOR2XL U11406 ( .A(n18776), .B(n18773), .Y(n13020) );
  NOR2XL U11407 ( .A(n18780), .B(n18779), .Y(n13019) );
  NAND4XL U11408 ( .A(n18776), .B(n18773), .C(n18780), .D(n18779), .Y(n13001)
         );
  NAND4XL U11409 ( .A(n18767), .B(n18770), .C(n18786), .D(n18783), .Y(n13002)
         );
  XOR2XL U11410 ( .A(n11592), .B(n13012), .Y(n11608) );
  CMPR32X1 U11411 ( .A(n18767), .B(n11604), .C(n11603), .CO(n24042), .S(n25791) );
  OAI21XL U11412 ( .A0(n20602), .A1(n3073), .B0(n20601), .Y(n20635) );
  NAND2XL U11413 ( .A(n20600), .B(n20599), .Y(n20601) );
  NAND3XL U11414 ( .A(n20596), .B(n20595), .C(n20576), .Y(n20600) );
  XOR2XL U11415 ( .A(n7395), .B(n7845), .Y(n7415) );
  INVXL U11416 ( .A(n19073), .Y(n19057) );
  INVX1 U11417 ( .A(n20321), .Y(n20326) );
  NOR2X1 U11418 ( .A(n5989), .B(n5934), .Y(n5933) );
  XOR2XL U11419 ( .A(n18761), .B(n19031), .Y(n18782) );
  NOR2XL U11420 ( .A(n15849), .B(n3077), .Y(n15850) );
  NOR2XL U11421 ( .A(n21008), .B(n15688), .Y(n15842) );
  NOR2XL U11422 ( .A(n15898), .B(n3077), .Y(n15855) );
  NOR2XL U11423 ( .A(n25006), .B(n15688), .Y(n15880) );
  NOR2XL U11424 ( .A(n21007), .B(n21006), .Y(n21011) );
  NOR2XL U11425 ( .A(n22266), .B(n22124), .Y(n22270) );
  NAND2XL U11426 ( .A(n23350), .B(n23316), .Y(n22378) );
  INVXL U11427 ( .A(n22271), .Y(n22315) );
  NAND2XL U11428 ( .A(n22313), .B(n22312), .Y(n22314) );
  INVX2 U11429 ( .A(n5569), .Y(n23864) );
  NOR2X2 U11430 ( .A(n7871), .B(n5603), .Y(n23863) );
  NOR2X1 U11431 ( .A(n7878), .B(n23199), .Y(n5603) );
  NOR2XL U11432 ( .A(n10720), .B(n7877), .Y(n7878) );
  NAND3X1 U11433 ( .A(n4671), .B(n3894), .C(n3895), .Y(n20673) );
  XOR2X1 U11434 ( .A(M3_mult_x_15_b_1_), .B(n18118), .Y(n6038) );
  XNOR2X1 U11435 ( .A(n21054), .B(n25876), .Y(n6362) );
  XNOR2X1 U11436 ( .A(n12265), .B(M3_mult_x_15_b_1_), .Y(n12266) );
  OAI22XL U11437 ( .A0(n18177), .A1(M3_mult_x_15_b_1_), .B0(n18165), .B1(
        n18223), .Y(n18161) );
  INVXL U11438 ( .A(n8569), .Y(n8247) );
  INVXL U11439 ( .A(n19641), .Y(n19448) );
  INVXL U11440 ( .A(n19663), .Y(n19377) );
  NAND2XL U11441 ( .A(n21643), .B(n21674), .Y(n21536) );
  INVXL U11442 ( .A(n21671), .Y(n21543) );
  NAND2XL U11443 ( .A(n21689), .B(n21708), .Y(n21542) );
  INVXL U11444 ( .A(n21678), .Y(n21546) );
  NAND2XL U11445 ( .A(n21689), .B(n21544), .Y(n21545) );
  NAND2XL U11446 ( .A(n21580), .B(n21563), .Y(n21477) );
  INVXL U11447 ( .A(n21708), .Y(n21523) );
  NAND2XL U11448 ( .A(n21643), .B(n21678), .Y(n21522) );
  OAI22XL U11449 ( .A0(n7511), .A1(n7051), .B0(n7512), .B1(n7050), .Y(n7054)
         );
  NAND2BXL U11450 ( .AN(n6944), .B(n25867), .Y(n6606) );
  XNOR2XL U11451 ( .A(n4806), .B(n3209), .Y(n6615) );
  XNOR2XL U11452 ( .A(n4806), .B(n25869), .Y(n6327) );
  XNOR2X2 U11453 ( .A(n6476), .B(M0_a_12_), .Y(n6298) );
  XNOR2XL U11454 ( .A(n16614), .B(M3_mult_x_15_b_1_), .Y(n16615) );
  XNOR2XL U11455 ( .A(n3203), .B(n11499), .Y(n16468) );
  XOR2X1 U11456 ( .A(M5_mult_x_15_n1), .B(n5718), .Y(n16108) );
  XNOR2XL U11457 ( .A(n5677), .B(M3_mult_x_15_b_1_), .Y(n16374) );
  XNOR2XL U11458 ( .A(n23221), .B(n25877), .Y(n7232) );
  NOR2X1 U11459 ( .A(n25243), .B(n23991), .Y(n5492) );
  INVXL U11460 ( .A(n9966), .Y(n6062) );
  OAI22XL U11461 ( .A0(n12597), .A1(n12201), .B0(n12595), .B1(n12171), .Y(
        n12188) );
  OAI22XL U11462 ( .A0(n13085), .A1(n13721), .B0(n13115), .B1(n13790), .Y(
        n13095) );
  NAND2BXL U11463 ( .AN(n13049), .B(n13898), .Y(n13084) );
  XNOR2X1 U11464 ( .A(n13769), .B(n13844), .Y(n13094) );
  NAND2X2 U11465 ( .A(n25229), .B(target_temp[11]), .Y(n6049) );
  CLKINVX3 U11466 ( .A(n13842), .Y(n13844) );
  OAI22XL U11467 ( .A0(n18624), .A1(n18603), .B0(n18625), .B1(n17905), .Y(
        n17908) );
  NAND2BXL U11468 ( .AN(n2978), .B(n18604), .Y(n17905) );
  OAI22X1 U11469 ( .A0(n17904), .A1(n18223), .B0(n18226), .B1(n17934), .Y(
        n4882) );
  OAI22XL U11470 ( .A0(n18239), .A1(n18142), .B0(n18141), .B1(n18140), .Y(
        n18153) );
  XNOR2XL U11471 ( .A(n18150), .B(n11499), .Y(n18104) );
  XNOR2XL U11472 ( .A(n3206), .B(n3197), .Y(n18241) );
  NAND2BXL U11473 ( .AN(n2978), .B(n18468), .Y(n17964) );
  XOR2X1 U11474 ( .A(M3_mult_x_15_b_1_), .B(n3210), .Y(n6129) );
  OAI21XL U11475 ( .A0(n25243), .A1(n25911), .B0(n11535), .Y(M1_a_16_) );
  OAI21XL U11476 ( .A0(n25243), .A1(n25910), .B0(n11539), .Y(M1_a_17_) );
  INVXL U11477 ( .A(n23204), .Y(n19411) );
  INVXL U11478 ( .A(n23205), .Y(n19404) );
  AOI2BB2XL U11479 ( .B0(n15190), .B1(n14987), .A0N(n15558), .A1N(n15436), .Y(
        n15302) );
  XNOR2XL U11480 ( .A(n23221), .B(n25876), .Y(n7290) );
  AOI222XL U11481 ( .A0(n22932), .A1(n23109), .B0(n22904), .B1(n11062), .C0(
        n22931), .C1(n3217), .Y(n22933) );
  XOR2XL U11482 ( .A(n22918), .B(n3056), .Y(M6_mult_x_15_n1105) );
  INVXL U11483 ( .A(n10811), .Y(n10824) );
  CMPR32X1 U11484 ( .A(n6455), .B(n6454), .C(n6453), .CO(n6467), .S(n6701) );
  ADDFX2 U11485 ( .A(n6484), .B(n6483), .CI(n6482), .CO(n6533), .S(n6505) );
  OAI22XL U11486 ( .A0(n7511), .A1(n6476), .B0(n7512), .B1(n6475), .Y(n6483)
         );
  NAND2BXL U11487 ( .AN(n6944), .B(n25868), .Y(n6475) );
  ADDFX2 U11488 ( .A(n6527), .B(n6526), .CI(n6525), .CO(n6689), .S(n6543) );
  NOR2BXL U11489 ( .AN(n6944), .B(n7556), .Y(n6527) );
  OAI22XL U11490 ( .A0(n6845), .A1(n6471), .B0(n6470), .B1(n6843), .Y(n6526)
         );
  XNOR2XL U11491 ( .A(n4806), .B(n23221), .Y(n6348) );
  AOI22XL U11492 ( .A0(n6733), .A1(target_temp[13]), .B0(n3229), .B1(w1[13]), 
        .Y(n6265) );
  XNOR2XL U11493 ( .A(n10858), .B(n10857), .Y(n22924) );
  NAND2XL U11494 ( .A(n10856), .B(n10855), .Y(n10857) );
  AOI21XL U11495 ( .A0(n10853), .A1(n10852), .B0(n10851), .Y(n10858) );
  INVXL U11496 ( .A(n10854), .Y(n10856) );
  NOR2BXL U11497 ( .AN(n3110), .B(n3105), .Y(n16530) );
  OAI22X1 U11498 ( .A0(n16638), .A1(n16396), .B0(n16341), .B1(n16475), .Y(
        n16399) );
  NOR2BXL U11499 ( .AN(n3110), .B(n17061), .Y(n16400) );
  CMPR32X1 U11500 ( .A(n16414), .B(n16413), .C(n16412), .CO(n16458), .S(n16484) );
  OAI22XL U11501 ( .A0(n16701), .A1(n16459), .B0(n16699), .B1(n16345), .Y(
        n16414) );
  XNOR2XL U11502 ( .A(n3203), .B(M3_mult_x_15_b_9_), .Y(n16373) );
  XNOR2XL U11503 ( .A(n3211), .B(n2974), .Y(n16382) );
  XNOR2XL U11504 ( .A(n5677), .B(M3_mult_x_15_b_2_), .Y(n16072) );
  CMPR32X1 U11505 ( .A(n9365), .B(n9364), .C(n9363), .CO(n9471), .S(n9334) );
  AOI22X1 U11506 ( .A0(n9164), .A1(y12[15]), .B0(n14427), .B1(y10[15]), .Y(
        n9046) );
  AOI22X1 U11507 ( .A0(n4566), .A1(data[21]), .B0(in_valid_d), .B1(w1[277]), 
        .Y(n9064) );
  NOR2BXL U11508 ( .AN(n9960), .B(n10403), .Y(n9752) );
  OAI22X1 U11509 ( .A0(n9782), .A1(n3180), .B0(n9963), .B1(n5296), .Y(n9801)
         );
  NOR2BXL U11510 ( .AN(n9960), .B(n9780), .Y(n9802) );
  NAND2BXL U11511 ( .AN(n9960), .B(n10324), .Y(n9799) );
  XNOR2X1 U11512 ( .A(n10324), .B(n10311), .Y(n9600) );
  NAND2X1 U11513 ( .A(n11536), .B(n4724), .Y(n5251) );
  NAND2X1 U11514 ( .A(n14427), .B(y10[12]), .Y(n5253) );
  NAND2X1 U11515 ( .A(n4856), .B(y12[12]), .Y(n5252) );
  NOR2X1 U11516 ( .A(n25243), .B(n23990), .Y(n5505) );
  OAI211X1 U11517 ( .A0(n23988), .A1(n25243), .B0(n9067), .C0(n11537), .Y(
        M2_b_18_) );
  XOR2X1 U11518 ( .A(M2_a_7_), .B(M2_a_6_), .Y(n5343) );
  XNOR2X1 U11519 ( .A(n12282), .B(n12560), .Y(n12105) );
  XNOR2XL U11520 ( .A(n14266), .B(M1_b_19_), .Y(n14079) );
  XOR2XL U11521 ( .A(n5430), .B(n3210), .Y(n5769) );
  XNOR2X1 U11522 ( .A(n18500), .B(M3_mult_x_15_b_9_), .Y(n17870) );
  BUFX3 U11523 ( .A(n18226), .Y(n18177) );
  BUFX3 U11524 ( .A(M1_a_2_), .Y(n13864) );
  BUFX3 U11525 ( .A(M1_a_6_), .Y(n14028) );
  NOR2XL U11526 ( .A(n14228), .B(n5391), .Y(M1_U4_U1_enc_tree_1__1__14_) );
  BUFX1 U11527 ( .A(n14119), .Y(n5512) );
  NOR2XL U11528 ( .A(n4807), .B(n4848), .Y(M1_U4_U1_or2_tree_0__1__24_) );
  OAI21XL U11529 ( .A0(n25243), .A1(n25904), .B0(n11517), .Y(M1_a_8_) );
  OAI21XL U11530 ( .A0(n25243), .A1(n25908), .B0(n11532), .Y(M1_a_15_) );
  OAI21XL U11531 ( .A0(n25243), .A1(n26235), .B0(n11525), .Y(M1_a_13_) );
  XNOR2XL U11532 ( .A(n14357), .B(n25861), .Y(n14057) );
  NAND2X2 U11533 ( .A(n25229), .B(target_temp[15]), .Y(n11527) );
  BUFX3 U11534 ( .A(M1_a_12_), .Y(n14196) );
  XOR2XL U11535 ( .A(n4164), .B(n3198), .Y(n5760) );
  CLKINVX3 U11536 ( .A(M1_b_15_), .Y(n14197) );
  XNOR2XL U11537 ( .A(n14266), .B(n14030), .Y(n13699) );
  OAI22X1 U11538 ( .A0(n13723), .A1(n14291), .B0(n13696), .B1(n6191), .Y(
        n13732) );
  OAI21X2 U11539 ( .A0(n13714), .A1(n3173), .B0(n6054), .Y(n6053) );
  NAND2X1 U11540 ( .A(n6056), .B(n6055), .Y(n6054) );
  OR2XL U11541 ( .A(n8456), .B(n8614), .Y(n8458) );
  AOI21XL U11542 ( .A0(n8442), .A1(n8823), .B0(n3155), .Y(n8441) );
  AOI22XL U11543 ( .A0(n8439), .A1(n8438), .B0(n8785), .B1(n8610), .Y(n8440)
         );
  OAI21XL U11544 ( .A0(n3160), .A1(n8400), .B0(n8399), .Y(n8641) );
  AOI21XL U11545 ( .A0(n8400), .A1(n8823), .B0(n3155), .Y(n8399) );
  OAI21XL U11546 ( .A0(n8398), .A1(n8397), .B0(n8493), .Y(n8400) );
  AOI22XL U11547 ( .A0(n19716), .A1(n19715), .B0(n19914), .B1(n19730), .Y(
        n19717) );
  OR2XL U11548 ( .A(n19733), .B(n19748), .Y(n19735) );
  OAI21XL U11549 ( .A0(n3165), .A1(n19454), .B0(n19453), .Y(n19775) );
  AOI21XL U11550 ( .A0(n19454), .A1(n19952), .B0(n3164), .Y(n19453) );
  OAI211XL U11551 ( .A0(n19807), .A1(n19576), .B0(n19424), .C0(n19452), .Y(
        n19454) );
  NAND2XL U11552 ( .A(n19553), .B(n19807), .Y(n19452) );
  NAND2XL U11553 ( .A(n15190), .B(n15006), .Y(n15007) );
  NAND2XL U11554 ( .A(n15190), .B(n14989), .Y(n14990) );
  AOI2BB2XL U11555 ( .B0(n15008), .B1(n15228), .A0N(n15008), .A1N(n15260), .Y(
        n15306) );
  AOI2BB2XL U11556 ( .B0(n15008), .B1(n15226), .A0N(n15008), .A1N(n15243), .Y(
        n15305) );
  AOI2BB2XL U11557 ( .B0(n15558), .B1(n14998), .A0N(n15558), .A1N(n15098), .Y(
        n15304) );
  NOR2XL U11558 ( .A(n15289), .B(n15305), .Y(n15352) );
  NAND2XL U11559 ( .A(n15019), .B(n15022), .Y(n15020) );
  AOI22XL U11560 ( .A0(n3095), .A1(n21564), .B0(n21572), .B1(n21580), .Y(
        n21855) );
  AOI2BB2XL U11561 ( .B0(n3172), .B1(n21781), .A0N(n3172), .A1N(n21782), .Y(
        n21741) );
  AOI2BB2XL U11562 ( .B0(n3172), .B1(n21777), .A0N(n3172), .A1N(n21780), .Y(
        n21751) );
  OAI21XL U11563 ( .A0(n3160), .A1(n8377), .B0(n8376), .Y(n8639) );
  AOI21XL U11564 ( .A0(n8377), .A1(n8823), .B0(n3155), .Y(n8376) );
  AOI22XL U11565 ( .A0(n8374), .A1(n8373), .B0(n8610), .B1(n8805), .Y(n8375)
         );
  OAI21XL U11566 ( .A0(n3160), .A1(n8419), .B0(n8418), .Y(n8637) );
  AOI21XL U11567 ( .A0(n8419), .A1(n8823), .B0(n3155), .Y(n8418) );
  OAI21XL U11568 ( .A0(n8800), .A1(n8593), .B0(n8416), .Y(n8417) );
  NAND4XL U11569 ( .A(n7905), .B(n7904), .C(n7903), .D(n7902), .Y(n8480) );
  NAND2XL U11570 ( .A(n19346), .B(w2[1]), .Y(n7904) );
  NAND2XL U11571 ( .A(n6217), .B(y10[1]), .Y(n7905) );
  AOI222XL U11572 ( .A0(n23152), .A1(n11059), .B0(n23093), .B1(n11058), .C0(
        n23150), .C1(n23151), .Y(n23138) );
  AOI222XL U11573 ( .A0(n23152), .A1(n23151), .B0(n23093), .B1(n10789), .C0(
        n23150), .C1(n3220), .Y(n23153) );
  AOI222XL U11574 ( .A0(n22932), .A1(n11073), .B0(n22904), .B1(n11063), .C0(
        n22931), .C1(n23109), .Y(n22872) );
  XOR2XL U11575 ( .A(n22848), .B(n3056), .Y(M6_mult_x_15_n1101) );
  XOR2XL U11576 ( .A(n22938), .B(n3055), .Y(M6_mult_x_15_n1125) );
  NAND2XL U11577 ( .A(n23152), .B(n22987), .Y(n4707) );
  XOR2XL U11578 ( .A(n22762), .B(n22606), .Y(n23139) );
  NAND2XL U11579 ( .A(n22761), .B(n22759), .Y(n22606) );
  XOR2XL U11580 ( .A(n22570), .B(n22569), .Y(n23104) );
  NAND2XL U11581 ( .A(n22568), .B(n22567), .Y(n22569) );
  OAI21XL U11582 ( .A0(n6699), .A1(n6698), .B0(n6697), .Y(n5624) );
  NAND2BX1 U11583 ( .AN(n6669), .B(n5554), .Y(n5553) );
  OAI22XL U11584 ( .A0(n6991), .A1(n6302), .B0(n6990), .B1(n6286), .Y(n6306)
         );
  OAI22XL U11585 ( .A0(n7535), .A1(n6301), .B0(n6312), .B1(n7460), .Y(n6307)
         );
  NAND2BXL U11586 ( .AN(M0_b_1_), .B(n5578), .Y(n5577) );
  INVXL U11587 ( .A(n5577), .Y(M0_U4_U1_or2_tree_0__1__28_) );
  NAND2X1 U11588 ( .A(n6245), .B(n5584), .Y(M0_a_6_) );
  OAI21X2 U11589 ( .A0(n7382), .A1(n26015), .B0(n6239), .Y(M0_a_18_) );
  AOI21X1 U11590 ( .A0(n7389), .A1(y10[18]), .B0(n4771), .Y(n6239) );
  NOR2XL U11591 ( .A(n25867), .B(n3209), .Y(M0_U3_U1_or2_tree_0__1__24_) );
  NOR2X1 U11592 ( .A(n17167), .B(n26013), .Y(n5943) );
  NOR2XL U11593 ( .A(M3_a_11_), .B(M3_a_9_), .Y(M3_U3_U1_or2_tree_0__1__20_)
         );
  AOI21XL U11594 ( .A0(n22931), .A1(n3218), .B0(n22905), .Y(n22906) );
  OAI2BB1XL U11595 ( .A0N(n11071), .A1N(n22904), .B0(n22903), .Y(n22905) );
  XOR2XL U11596 ( .A(n10792), .B(n10791), .Y(n23148) );
  NAND2XL U11597 ( .A(n10790), .B(n11050), .Y(n10791) );
  INVXL U11598 ( .A(n11046), .Y(n10790) );
  INVXL U11599 ( .A(n22945), .Y(n22951) );
  AOI222XL U11600 ( .A0(n23152), .A1(n10769), .B0(n23093), .B1(n23002), .C0(
        n23150), .C1(n10749), .Y(n22944) );
  NAND2X1 U11601 ( .A(n16395), .B(n16394), .Y(n5702) );
  OR2X2 U11602 ( .A(n16395), .B(n16394), .Y(n5703) );
  OAI22X2 U11603 ( .A0(n15942), .A1(n26018), .B0(n25920), .B1(n15940), .Y(
        n5651) );
  NOR2XL U11604 ( .A(M4_a_13_), .B(M4_a_12_), .Y(M4_U3_U1_enc_tree_1__1__18_)
         );
  NOR2XL U11605 ( .A(M4_a_5_), .B(M4_a_4_), .Y(M4_U3_U1_enc_tree_1__1__26_) );
  NOR2XL U11606 ( .A(n18006), .B(M4_a_0_), .Y(M4_U3_U1_enc_tree_1__1__30_) );
  OAI22XL U11607 ( .A0(n10517), .A1(n9581), .B0(n10533), .B1(n10162), .Y(
        n10163) );
  INVXL U11608 ( .A(n9288), .Y(n4818) );
  XOR2X1 U11609 ( .A(n9248), .B(n5245), .Y(n5244) );
  OAI22XL U11610 ( .A0(n12535), .A1(M3_mult_x_15_b_3_), .B0(n12995), .B1(
        n11499), .Y(n11696) );
  XNOR2X1 U11611 ( .A(n12758), .B(n12271), .Y(n11728) );
  XNOR2XL U11612 ( .A(n2980), .B(n3202), .Y(n11727) );
  NAND2XL U11613 ( .A(n5779), .B(n12020), .Y(n5778) );
  XNOR2X1 U11614 ( .A(n12758), .B(M3_mult_x_15_b_1_), .Y(n11812) );
  XNOR2XL U11615 ( .A(n12732), .B(n3201), .Y(n12514) );
  CLKINVX3 U11616 ( .A(n4919), .Y(n4918) );
  OAI22XL U11617 ( .A0(n18111), .A1(n17903), .B0(n18504), .B1(n17893), .Y(
        n17888) );
  OAI21X1 U11618 ( .A0(n18239), .A1(n5815), .B0(n5814), .Y(n17887) );
  XNOR2X1 U11619 ( .A(n18503), .B(n18611), .Y(n17602) );
  INVX1 U11620 ( .A(M1_b_12_), .Y(n5488) );
  AOI21XL U11621 ( .A0(n3019), .A1(M1_b_18_), .B0(n5391), .Y(
        M1_U4_U1_enc_tree_0__1__14_) );
  XNOR2XL U11622 ( .A(n12732), .B(n3190), .Y(n11918) );
  OAI22X1 U11623 ( .A0(n17148), .A1(n3110), .B0(M3_mult_x_15_b_1_), .B1(n17147), .Y(n15974) );
  OAI21XL U11624 ( .A0(n3194), .A1(n3110), .B0(n17148), .Y(n15975) );
  OAI22X2 U11625 ( .A0(n18522), .A1(n17518), .B0(n17509), .B1(n3195), .Y(n5864) );
  XNOR2X1 U11626 ( .A(n18453), .B(n12561), .Y(n17552) );
  OAI22XL U11627 ( .A0(n18522), .A1(n17582), .B0(n3195), .B1(n17518), .Y(
        n17549) );
  OAI2BB1X1 U11628 ( .A0N(n13665), .A1N(n13664), .B0(n13663), .Y(n13706) );
  NAND2XL U11629 ( .A(n8641), .B(n8640), .Y(n8931) );
  AOI21XL U11630 ( .A0(n19809), .A1(n19952), .B0(n3164), .Y(n19808) );
  OAI211XL U11631 ( .A0(n19807), .A1(n19806), .B0(n19424), .C0(n19805), .Y(
        n19809) );
  AOI21XL U11632 ( .A0(n19801), .A1(n19952), .B0(n3164), .Y(n19800) );
  OAI211XL U11633 ( .A0(n19807), .A1(n19799), .B0(n19424), .C0(n19798), .Y(
        n19801) );
  NOR2XL U11634 ( .A(n19981), .B(n19985), .Y(n19988) );
  INVXL U11635 ( .A(n19980), .Y(n19981) );
  INVXL U11636 ( .A(n19910), .Y(n19989) );
  AOI21XL U11637 ( .A0(n19840), .A1(n19952), .B0(n3164), .Y(n19839) );
  NAND2XL U11638 ( .A(n19424), .B(n19838), .Y(n19840) );
  INVXL U11639 ( .A(n20060), .Y(n19770) );
  INVXL U11640 ( .A(n20054), .Y(n19771) );
  NOR2XL U11641 ( .A(n23210), .B(n23209), .Y(n19342) );
  NOR2XL U11642 ( .A(n23206), .B(n23205), .Y(n19344) );
  OAI211XL U11643 ( .A0(n3090), .A1(n15419), .B0(n15046), .C0(n15418), .Y(
        n15421) );
  NAND2XL U11644 ( .A(n22131), .B(n22130), .Y(n22093) );
  NOR2X1 U11645 ( .A(n23406), .B(n21446), .Y(n21481) );
  NAND2XL U11646 ( .A(n21331), .B(w1[21]), .Y(n21308) );
  NAND2XL U11647 ( .A(n21311), .B(temp0[0]), .Y(n21190) );
  NAND2XL U11648 ( .A(n21256), .B(temp0[4]), .Y(n21174) );
  NAND2XL U11649 ( .A(n21329), .B(temp0[14]), .Y(n21255) );
  NAND2XL U11650 ( .A(n21333), .B(temp0[15]), .Y(n21250) );
  INVXL U11651 ( .A(n21517), .Y(n21978) );
  NAND2BXL U11652 ( .AN(n21712), .B(n21507), .Y(n21742) );
  OAI22X1 U11653 ( .A0(n11642), .A1(n12635), .B0(n12633), .B1(n6040), .Y(
        n11780) );
  INVXL U11654 ( .A(n11694), .Y(n4955) );
  XNOR2XL U11655 ( .A(M3_mult_x_15_b_20_), .B(n3211), .Y(n5947) );
  XOR2XL U11656 ( .A(n22883), .B(n3119), .Y(M6_mult_x_15_n1044) );
  XOR2XL U11657 ( .A(n22914), .B(n3053), .Y(M6_mult_x_15_n1164) );
  XOR2XL U11658 ( .A(n22670), .B(n3055), .Y(M6_mult_x_15_n1116) );
  XOR2XL U11659 ( .A(n22910), .B(n3058), .Y(M6_mult_x_15_n1068) );
  XOR2XL U11660 ( .A(n22936), .B(n3056), .Y(M6_mult_x_15_n1092) );
  XOR2XL U11661 ( .A(n22877), .B(n3119), .Y(M6_mult_x_15_n1048) );
  XOR2XL U11662 ( .A(n22879), .B(n3058), .Y(M6_mult_x_15_n1072) );
  XOR2XL U11663 ( .A(n22965), .B(n3055), .Y(M6_mult_x_15_n1120) );
  XOR2XL U11664 ( .A(n22529), .B(n22501), .Y(n22800) );
  NAND2XL U11665 ( .A(n22528), .B(n22526), .Y(n22501) );
  AOI222XL U11666 ( .A0(n22932), .A1(n9109), .B0(n22904), .B1(n11074), .C0(
        n22931), .C1(n3219), .Y(n22810) );
  NAND2X1 U11667 ( .A(n5604), .B(w2[21]), .Y(n5605) );
  NAND2X1 U11668 ( .A(n6733), .B(y10[21]), .Y(n5606) );
  OAI22X1 U11669 ( .A0(n18522), .A1(n17508), .B0(n3195), .B1(n17636), .Y(
        n17618) );
  XOR2XL U11670 ( .A(n22682), .B(n3221), .Y(M6_mult_x_15_n1192) );
  XOR2XL U11671 ( .A(n22731), .B(n3053), .Y(M6_mult_x_15_n1168) );
  XOR2XL U11672 ( .A(n22852), .B(n3054), .Y(M6_mult_x_15_n1144) );
  OAI22X2 U11673 ( .A0(n15942), .A1(n26031), .B0(n26271), .B1(n15940), .Y(
        n4941) );
  INVX1 U11674 ( .A(M5_a_4_), .Y(n4783) );
  OAI222X1 U11675 ( .A0(n26041), .A1(n15941), .B0(n25933), .B1(n25813), .C0(
        n26281), .C1(n15940), .Y(M5_a_4_) );
  NAND3X2 U11676 ( .A(n5728), .B(n5727), .C(n5726), .Y(M5_a_8_) );
  NAND2XL U11677 ( .A(n4875), .B(data[104]), .Y(n5727) );
  OAI22X2 U11678 ( .A0(n4860), .A1(n26019), .B0(n25921), .B1(n17167), .Y(n5639) );
  NOR2X1 U11679 ( .A(n4860), .B(n26446), .Y(n5031) );
  OAI22X1 U11680 ( .A0(n17060), .A1(n5640), .B0(n15960), .B1(n17061), .Y(
        n16029) );
  ADDFX2 U11681 ( .A(n16034), .B(n16033), .CI(n16032), .CO(n16120), .S(n16038)
         );
  OAI22XL U11682 ( .A0(n16704), .A1(n15956), .B0(n5835), .B1(n3047), .Y(n16033) );
  NOR2XL U11683 ( .A(n23181), .B(n23180), .Y(n8214) );
  XOR2X1 U11684 ( .A(n5142), .B(n9716), .Y(n9763) );
  OAI22X1 U11685 ( .A0(n12152), .A1(n11634), .B0(n3185), .B1(n12265), .Y(
        n11760) );
  OAI22X1 U11686 ( .A0(n12618), .A1(n11640), .B0(n11781), .B1(n12616), .Y(
        n11761) );
  CMPR32X1 U11687 ( .A(n11774), .B(n11773), .C(n11772), .CO(n11875), .S(n11754) );
  OAI2BB1X1 U11688 ( .A0N(n11797), .A1N(n5787), .B0(n5785), .Y(n11804) );
  OAI21XL U11689 ( .A0(n4914), .A1(n4913), .B0(n4911), .Y(n12602) );
  INVXL U11690 ( .A(n12644), .Y(n4913) );
  NAND2XL U11691 ( .A(n4923), .B(n11834), .Y(n4922) );
  NAND2BXL U11692 ( .AN(n11835), .B(n4924), .Y(n4923) );
  CMPR32X1 U11693 ( .A(n3107), .B(n12580), .C(n12579), .CO(n12693), .S(n12569)
         );
  OAI22XL U11694 ( .A0(n12618), .A1(n25884), .B0(n12616), .B1(n3191), .Y(
        n12579) );
  OAI22XL U11695 ( .A0(n12535), .A1(n3198), .B0(n12995), .B1(n3021), .Y(n12580) );
  OAI22XL U11696 ( .A0(n18083), .A1(n17707), .B0(n18429), .B1(n17671), .Y(
        n17723) );
  NOR2BXL U11697 ( .AN(n13049), .B(n14356), .Y(n13599) );
  ADDFX2 U11698 ( .A(n17782), .B(n17781), .CI(n17780), .CO(n17819), .S(n17772)
         );
  OAI22X1 U11699 ( .A0(n18659), .A1(n17777), .B0(n17832), .B1(n17833), .Y(
        n17824) );
  CMPR32X1 U11700 ( .A(n12630), .B(n12629), .C(n12628), .CO(n12653), .S(n12649) );
  OAI22XL U11701 ( .A0(n12717), .A1(n11978), .B0(n12718), .B1(n12593), .Y(
        n12630) );
  CMPR32X1 U11702 ( .A(n11983), .B(n11982), .C(n11981), .CO(n12648), .S(n11970) );
  OAI22XL U11703 ( .A0(n12635), .A1(n11951), .B0(n12633), .B1(n11980), .Y(
        n11982) );
  OAI22XL U11704 ( .A0(n18541), .A1(n17654), .B0(n5893), .B1(n17535), .Y(
        n17664) );
  OAI21XL U11705 ( .A0(n17599), .A1(n17598), .B0(n17597), .Y(n5035) );
  INVXL U11706 ( .A(n14499), .Y(n14333) );
  NAND2X1 U11707 ( .A(n21166), .B(sigma11[21]), .Y(n6095) );
  AOI22XL U11708 ( .A0(n5480), .A1(sigma11[22]), .B0(in_valid_t), .B1(w2[54]), 
        .Y(n17478) );
  NOR2XL U11709 ( .A(n8852), .B(n8856), .Y(n8859) );
  INVXL U11710 ( .A(n8851), .Y(n8852) );
  NAND2XL U11711 ( .A(n8921), .B(n8920), .Y(n8922) );
  INVXL U11712 ( .A(n8919), .Y(n8921) );
  NAND2XL U11713 ( .A(n19829), .B(n19828), .Y(n19866) );
  NAND2XL U11714 ( .A(n19835), .B(n19834), .Y(n19853) );
  NAND2XL U11715 ( .A(n19825), .B(n19824), .Y(n19879) );
  NAND2XL U11716 ( .A(n19833), .B(n19832), .Y(n19857) );
  NAND2XL U11717 ( .A(n19827), .B(n19826), .Y(n19874) );
  INVXL U11718 ( .A(n20186), .Y(n20219) );
  NAND2XL U11719 ( .A(n21331), .B(w1[14]), .Y(n21254) );
  INVXL U11720 ( .A(n21514), .Y(n21962) );
  NAND2XL U11721 ( .A(n21333), .B(w1[19]), .Y(n21294) );
  NAND2XL U11722 ( .A(n21466), .B(n21480), .Y(n21467) );
  INVXL U11723 ( .A(n21478), .Y(n21466) );
  NAND2XL U11724 ( .A(n21311), .B(temp0[20]), .Y(n21293) );
  NAND2XL U11725 ( .A(n21331), .B(temp0[22]), .Y(n21312) );
  NAND2XL U11726 ( .A(n21256), .B(temp0[19]), .Y(n21295) );
  NAND2XL U11727 ( .A(n21329), .B(temp0[21]), .Y(n21309) );
  NAND2XL U11728 ( .A(n21329), .B(temp0[5]), .Y(n21216) );
  NOR2XL U11729 ( .A(n21224), .B(n21556), .Y(n21212) );
  OAI21XL U11730 ( .A0(n6193), .A1(n21256), .B0(n21241), .Y(n21473) );
  NAND2XL U11731 ( .A(n21331), .B(temp0[10]), .Y(n21241) );
  NAND2XL U11732 ( .A(n21311), .B(temp0[16]), .Y(n21248) );
  NAND2XL U11733 ( .A(n21333), .B(temp0[13]), .Y(n21253) );
  NAND2XL U11734 ( .A(n21331), .B(temp0[9]), .Y(n21242) );
  NOR2XL U11735 ( .A(n21265), .B(n21475), .Y(n21239) );
  NAND2XL U11736 ( .A(n15653), .B(n15652), .Y(n15654) );
  NAND2XL U11737 ( .A(n15682), .B(n15681), .Y(n15683) );
  NAND2XL U11738 ( .A(n15671), .B(n15670), .Y(n15672) );
  INVXL U11739 ( .A(n15669), .Y(n15671) );
  NAND2XL U11740 ( .A(n21885), .B(n21884), .Y(n21939) );
  NAND2XL U11741 ( .A(n21883), .B(n21882), .Y(n21944) );
  INVXL U11742 ( .A(n21970), .Y(n22048) );
  INVXL U11743 ( .A(n21963), .Y(n22041) );
  NOR2XL U11744 ( .A(n22040), .B(n22044), .Y(n22047) );
  INVXL U11745 ( .A(n22039), .Y(n22040) );
  NAND4XL U11746 ( .A(n19076), .B(n5602), .C(n20951), .D(n10738), .Y(n7319) );
  OAI2BB1XL U11747 ( .A0N(n6012), .A1N(n16964), .B0(n6011), .Y(n16988) );
  BUFX3 U11748 ( .A(n6828), .Y(n25872) );
  OAI2BB1XL U11749 ( .A0N(n5052), .A1N(n17091), .B0(n5051), .Y(n17098) );
  NAND2XL U11750 ( .A(n18840), .B(n13031), .Y(n12965) );
  NAND2X2 U11751 ( .A(n12494), .B(n12495), .Y(n12875) );
  NAND2XL U11752 ( .A(n18840), .B(n17414), .Y(n17288) );
  NOR2XL U11753 ( .A(M4_a_7_), .B(M4_a_5_), .Y(M4_U3_U1_or2_tree_0__1__24_) );
  INVXL U11754 ( .A(n7721), .Y(n7703) );
  ADDFX2 U11755 ( .A(n10524), .B(n10523), .CI(n10522), .CO(n10558), .S(n10552)
         );
  NAND2XL U11756 ( .A(n10558), .B(n10557), .Y(n10600) );
  INVXL U11757 ( .A(n10575), .Y(n10601) );
  NAND2XL U11758 ( .A(n10263), .B(n10262), .Y(n10277) );
  XOR2X1 U11759 ( .A(n17739), .B(n5887), .Y(n5886) );
  NOR2X2 U11760 ( .A(n18870), .B(n18881), .Y(n18419) );
  NAND2XL U11761 ( .A(n8746), .B(n8745), .Y(n8747) );
  INVXL U11762 ( .A(n8741), .Y(n8744) );
  NAND2XL U11763 ( .A(n8738), .B(n8737), .Y(n8739) );
  INVXL U11764 ( .A(n8736), .Y(n8738) );
  NAND2XL U11765 ( .A(n8725), .B(n8724), .Y(n8726) );
  INVXL U11766 ( .A(n8723), .Y(n8725) );
  NAND2XL U11767 ( .A(n8716), .B(n8855), .Y(n8717) );
  INVXL U11768 ( .A(n8856), .Y(n8716) );
  NAND2XL U11769 ( .A(n8729), .B(n8728), .Y(n8730) );
  NAND3XL U11770 ( .A(n20404), .B(n20457), .C(n20543), .Y(n9023) );
  OAI31XL U11771 ( .A0(n24798), .A1(n24716), .A2(n20112), .B0(n20111), .Y(
        n20113) );
  AOI211XL U11772 ( .A0(n20110), .A1(n20109), .B0(n24717), .C0(n24680), .Y(
        n20112) );
  AOI211XL U11773 ( .A0(n20105), .A1(n20104), .B0(n20195), .C0(n20196), .Y(
        n20108) );
  NAND2XL U11774 ( .A(n15505), .B(n15504), .Y(n15506) );
  INVXL U11775 ( .A(n15503), .Y(n15505) );
  NAND2XL U11776 ( .A(n15514), .B(n15513), .Y(n15515) );
  INVXL U11777 ( .A(n15512), .Y(n15514) );
  NAND2XL U11778 ( .A(n15500), .B(n15499), .Y(n15501) );
  INVXL U11779 ( .A(n15498), .Y(n15500) );
  NOR2X1 U11780 ( .A(n21496), .B(n21495), .Y(n21723) );
  NAND2XL U11781 ( .A(n21492), .B(n21497), .Y(n21494) );
  INVXL U11782 ( .A(n21702), .Y(n21722) );
  AOI2BB2XL U11783 ( .B0(n23116), .B1(n21901), .A0N(n21628), .A1N(n21902), .Y(
        n21728) );
  NOR2X1 U11784 ( .A(n3171), .B(n3096), .Y(n21793) );
  AOI2BB2XL U11785 ( .B0(n23116), .B1(n21862), .A0N(n21628), .A1N(n21863), .Y(
        n21731) );
  CLKINVX2 U11786 ( .A(n21803), .Y(n21801) );
  NAND2XL U11787 ( .A(n21497), .B(n21491), .Y(n21499) );
  INVXL U11788 ( .A(n23118), .Y(n21498) );
  NAND2XL U11789 ( .A(n15478), .B(n15477), .Y(n15479) );
  NAND2XL U11790 ( .A(n15599), .B(n15598), .Y(n15600) );
  INVXL U11791 ( .A(n15597), .Y(n15599) );
  INVX1 U11792 ( .A(n15532), .Y(n15613) );
  INVXL U11793 ( .A(n22285), .Y(n22241) );
  NAND2XL U11794 ( .A(n3126), .B(n22286), .Y(n22240) );
  NAND2XL U11795 ( .A(n3126), .B(n22282), .Y(n22255) );
  INVXL U11796 ( .A(n22282), .Y(n22283) );
  INVX1 U11797 ( .A(n21972), .Y(n22051) );
  AOI211XL U11798 ( .A0(n22160), .A1(n22159), .B0(n22286), .C0(n22287), .Y(
        n22162) );
  AOI211XL U11799 ( .A0(n22155), .A1(n22154), .B0(n22296), .C0(n22297), .Y(
        n22158) );
  NOR2X1 U11800 ( .A(n22448), .B(n22256), .Y(n22167) );
  NOR2XL U11801 ( .A(n22019), .B(n22023), .Y(n22014) );
  AOI21XL U11802 ( .A0(n7668), .A1(n7755), .B0(n7667), .Y(n7669) );
  NAND2XL U11803 ( .A(n7346), .B(n7345), .Y(n10732) );
  NAND2XL U11804 ( .A(n7347), .B(n7338), .Y(n7346) );
  AOI22XL U11805 ( .A0(n7344), .A1(n7343), .B0(n7342), .B1(n7341), .Y(n7345)
         );
  XOR2XL U11806 ( .A(n7337), .B(n7336), .Y(n7338) );
  NOR2XL U11807 ( .A(n7359), .B(n7358), .Y(n10734) );
  NAND2BXL U11808 ( .AN(n7357), .B(n7356), .Y(n7358) );
  INVXL U11809 ( .A(n7347), .Y(n7359) );
  XOR2XL U11810 ( .A(n7355), .B(n7354), .Y(n7356) );
  OAI21X1 U11811 ( .A0(n17388), .A1(n17391), .B0(n17392), .Y(n17362) );
  NOR2XL U11812 ( .A(n10946), .B(n10985), .Y(n10948) );
  NAND2XL U11813 ( .A(n10986), .B(n10944), .Y(n10946) );
  INVXL U11814 ( .A(n20542), .Y(n20545) );
  INVXL U11815 ( .A(n20562), .Y(n20397) );
  NAND2XL U11816 ( .A(n3067), .B(n20542), .Y(n20396) );
  NOR2XL U11817 ( .A(n3067), .B(n20580), .Y(n20401) );
  INVXL U11818 ( .A(n20402), .Y(n20403) );
  INVXL U11819 ( .A(n20561), .Y(n20564) );
  NAND2XL U11820 ( .A(n3067), .B(n20562), .Y(n20563) );
  INVXL U11821 ( .A(n20404), .Y(n20579) );
  NOR2X1 U11822 ( .A(n10618), .B(n10504), .Y(n10626) );
  INVXL U11823 ( .A(n15577), .Y(n15578) );
  INVXL U11824 ( .A(n15619), .Y(n15582) );
  NAND3XL U11825 ( .A(n25270), .B(n15860), .C(n21000), .Y(n15779) );
  NAND4XL U11826 ( .A(n15777), .B(n15923), .C(n15873), .D(n15920), .Y(n15778)
         );
  NAND2XL U11827 ( .A(n10663), .B(n10662), .Y(n10664) );
  AOI21XL U11828 ( .A0(n10277), .A1(n10265), .B0(n10264), .Y(n10706) );
  OAI22XL U11829 ( .A0(n10263), .A1(n10262), .B0(M2_U3_U1_enc_tree_4__4__16_), 
        .B1(n10261), .Y(n10264) );
  XOR2XL U11830 ( .A(n10259), .B(n10258), .Y(n10265) );
  INVXL U11831 ( .A(n10260), .Y(n10261) );
  NAND2XL U11832 ( .A(n10277), .B(n10276), .Y(n10708) );
  NOR2XL U11833 ( .A(n10275), .B(n10274), .Y(n10276) );
  XOR2XL U11834 ( .A(n10273), .B(n10272), .Y(n10274) );
  XNOR2XL U11835 ( .A(n10269), .B(n10268), .Y(n10275) );
  OAI21XL U11836 ( .A0(n14608), .A1(n14638), .B0(n14607), .Y(n14613) );
  INVXL U11837 ( .A(n14609), .Y(n14611) );
  INVXL U11838 ( .A(n14585), .Y(n14587) );
  AND4XL U11839 ( .A(n24285), .B(n25184), .C(n24087), .D(n24336), .Y(n11621)
         );
  INVXL U11840 ( .A(n19956), .Y(n19957) );
  NAND4XL U11841 ( .A(n24889), .B(n20255), .C(n24849), .D(n24717), .Y(n20165)
         );
  INVXL U11842 ( .A(n20235), .Y(n20238) );
  NAND2XL U11843 ( .A(n20001), .B(n20000), .Y(n20002) );
  INVXL U11844 ( .A(n19998), .Y(n19961) );
  NOR2XL U11845 ( .A(n23121), .B(n23120), .Y(n21441) );
  NOR2XL U11846 ( .A(n23125), .B(n23124), .Y(n21439) );
  NOR2XL U11847 ( .A(n21803), .B(n3171), .Y(n21702) );
  INVXL U11848 ( .A(n22287), .Y(n22243) );
  NAND2XL U11849 ( .A(n3126), .B(n22272), .Y(n22242) );
  AOI22X1 U11850 ( .A0(n22191), .A1(n22426), .B0(n22237), .B1(n3129), .Y(
        n22359) );
  INVXL U11851 ( .A(n22192), .Y(n22191) );
  INVXL U11852 ( .A(n22286), .Y(n22289) );
  NAND2XL U11853 ( .A(n3126), .B(n22287), .Y(n22288) );
  INVXL U11854 ( .A(n22272), .Y(n22275) );
  NAND2XL U11855 ( .A(n3126), .B(n22273), .Y(n22274) );
  AOI21XL U11856 ( .A0(n22344), .A1(n3129), .B0(n22300), .Y(n22373) );
  NOR2XL U11857 ( .A(n22341), .B(n3129), .Y(n22300) );
  NAND2XL U11858 ( .A(n3126), .B(n22333), .Y(n22253) );
  INVXL U11859 ( .A(n17383), .Y(n17385) );
  NAND4XL U11860 ( .A(n23468), .B(n19080), .C(n11466), .D(n11455), .Y(n11349)
         );
  NAND2XL U11861 ( .A(n4826), .B(target_temp[23]), .Y(n14455) );
  NAND2XL U11862 ( .A(n4826), .B(target_temp[26]), .Y(n14444) );
  NAND2XL U11863 ( .A(n4826), .B(target_temp[25]), .Y(n14448) );
  NOR2XL U11864 ( .A(n18767), .B(n18770), .Y(n13022) );
  INVXL U11865 ( .A(n20283), .Y(n23537) );
  NAND2XL U11866 ( .A(in_valid_t), .B(w2[27]), .Y(n11567) );
  NAND2XL U11867 ( .A(n21166), .B(sigma10[27]), .Y(n11568) );
  NAND2XL U11868 ( .A(n4875), .B(data[59]), .Y(n11569) );
  INVX1 U11869 ( .A(n19319), .Y(n19292) );
  NOR2X1 U11870 ( .A(n20284), .B(n20365), .Y(n5601) );
  NAND2XL U11871 ( .A(n10692), .B(n10676), .Y(n9189) );
  NAND2XL U11872 ( .A(n14600), .B(n14599), .Y(n14601) );
  INVXL U11873 ( .A(n14598), .Y(n14600) );
  INVXL U11874 ( .A(n14590), .Y(n14592) );
  OAI21XL U11875 ( .A0(n26302), .A1(n3115), .B0(n14414), .Y(n14704) );
  NAND2XL U11876 ( .A(in_valid_t), .B(w2[61]), .Y(n18756) );
  NAND2XL U11877 ( .A(n5032), .B(data[93]), .Y(n18758) );
  NAND2XL U11878 ( .A(n20232), .B(n20182), .Y(n20209) );
  INVXL U11879 ( .A(n20170), .Y(n20171) );
  NOR2XL U11880 ( .A(n22308), .B(n22307), .Y(n22309) );
  INVXL U11881 ( .A(n22305), .Y(n22306) );
  NAND2XL U11882 ( .A(n22237), .B(n22426), .Y(n22238) );
  NAND2X1 U11883 ( .A(n21336), .B(n21388), .Y(n21391) );
  AOI2BB2XL U11884 ( .B0(n22373), .B1(n3079), .A0N(n22372), .A1N(n3079), .Y(
        n22384) );
  NAND2XL U11885 ( .A(n23285), .B(n23297), .Y(n23261) );
  NAND2XL U11886 ( .A(n22362), .B(n3079), .Y(n22321) );
  AOI2BB2XL U11887 ( .B0(n22368), .B1(n3079), .A0N(n22367), .A1N(n3079), .Y(
        n22414) );
  NAND2XL U11888 ( .A(n22394), .B(n3082), .Y(n22435) );
  NAND2XL U11889 ( .A(n22393), .B(n3082), .Y(n22446) );
  NAND2XL U11890 ( .A(n23376), .B(n23380), .Y(n23369) );
  OAI21XL U11891 ( .A0(n6171), .A1(n21333), .B0(n21319), .Y(n21405) );
  NAND2XL U11892 ( .A(n21329), .B(temp0[27]), .Y(n21319) );
  NAND2XL U11893 ( .A(in_valid_t), .B(w2[57]), .Y(n18744) );
  NAND2XL U11894 ( .A(n3111), .B(data[89]), .Y(n18746) );
  NOR2XL U11895 ( .A(n7382), .B(n26042), .Y(n7374) );
  OAI2BB1XL U11896 ( .A0N(y10[24]), .A1N(n3224), .B0(n7400), .Y(n7859) );
  AOI22XL U11897 ( .A0(n6733), .A1(target_temp[24]), .B0(in_valid_d), .B1(
        w1[24]), .Y(n7400) );
  AOI22XL U11898 ( .A0(n7389), .A1(target_temp[30]), .B0(in_valid_d), .B1(
        w1[30]), .Y(n7369) );
  AOI22XL U11899 ( .A0(n6733), .A1(target_temp[23]), .B0(in_valid_d), .B1(
        w1[23]), .Y(n7401) );
  AOI22XL U11900 ( .A0(n6733), .A1(target_temp[25]), .B0(in_valid_d), .B1(
        w1[25]), .Y(n7398) );
  NOR2XL U11901 ( .A(n7382), .B(n26037), .Y(n7370) );
  NOR2XL U11902 ( .A(n7382), .B(n26036), .Y(n7372) );
  NAND2XL U11903 ( .A(in_valid_d), .B(w1[157]), .Y(n14430) );
  NAND2XL U11904 ( .A(n25233), .B(learning_rate[29]), .Y(n14431) );
  NAND4XL U11905 ( .A(n14456), .B(n14448), .C(n14447), .D(n14446), .Y(n14711)
         );
  NAND2XL U11906 ( .A(in_valid_d), .B(w1[153]), .Y(n14446) );
  NAND2XL U11907 ( .A(n25233), .B(learning_rate[25]), .Y(n14447) );
  AOI21XL U11908 ( .A0(n3223), .A1(sigma10[25]), .B0(n14409), .Y(n14701) );
  XOR2XL U11909 ( .A(n20823), .B(n20822), .Y(n23544) );
  NAND2XL U11910 ( .A(n23915), .B(n20821), .Y(n20823) );
  INVXL U11911 ( .A(n20820), .Y(n20821) );
  XOR2XL U11912 ( .A(n20299), .B(n20298), .Y(n23940) );
  NAND2XL U11913 ( .A(n23915), .B(n20297), .Y(n20299) );
  INVXL U11914 ( .A(n20296), .Y(n20297) );
  OR2XL U11915 ( .A(n20548), .B(n20547), .Y(n20549) );
  XOR2XL U11916 ( .A(n9142), .B(n10681), .Y(n9183) );
  INVXL U11917 ( .A(n20841), .Y(n24707) );
  NAND4XL U11918 ( .A(n23235), .B(n22229), .C(n22228), .D(n22227), .Y(n22230)
         );
  INVX1 U11919 ( .A(n23129), .Y(n22229) );
  NOR2XL U11920 ( .A(n20525), .B(n20576), .Y(n20514) );
  NOR2XL U11921 ( .A(n20502), .B(n20576), .Y(n20503) );
  NOR2XL U11922 ( .A(n20550), .B(n20597), .Y(n20498) );
  OAI22X1 U11923 ( .A0(n20540), .A1(n20539), .B0(n20538), .B1(n3073), .Y(
        n23754) );
  NOR2XL U11924 ( .A(n20577), .B(n20597), .Y(n20480) );
  XOR2XL U11925 ( .A(n7393), .B(n7847), .Y(n7413) );
  NAND2X1 U11926 ( .A(n3132), .B(n23492), .Y(n10712) );
  XOR2X2 U11927 ( .A(n19099), .B(n5190), .Y(n23521) );
  NOR2X1 U11928 ( .A(n20810), .B(n20707), .Y(n17489) );
  NOR2X1 U11929 ( .A(n20612), .B(n20810), .Y(n20613) );
  AND2X1 U11930 ( .A(n9188), .B(n9189), .Y(n20790) );
  XOR2X1 U11931 ( .A(n20986), .B(n20985), .Y(n23627) );
  NAND2X1 U11932 ( .A(n23744), .B(n20984), .Y(n20986) );
  INVXL U11933 ( .A(n20983), .Y(n20984) );
  NAND2X1 U11934 ( .A(n3134), .B(n5388), .Y(n5381) );
  XNOR2XL U11935 ( .A(n14700), .B(n14698), .Y(n14462) );
  XOR2XL U11936 ( .A(n14441), .B(n14705), .Y(n14468) );
  CMPR32X1 U11937 ( .A(n18767), .B(n18766), .C(n18765), .CO(n20651), .S(n25129) );
  NOR2XL U11938 ( .A(n24034), .B(n24033), .Y(n24037) );
  OR2XL U11939 ( .A(n24945), .B(n24944), .Y(n24946) );
  NOR2XL U11940 ( .A(n25280), .B(n15638), .Y(n24584) );
  NAND2XL U11941 ( .A(n15930), .B(n15929), .Y(n15931) );
  OAI22XL U11942 ( .A0(n24879), .A1(n24878), .B0(n3076), .B1(n24877), .Y(
        n24975) );
  NOR2XL U11943 ( .A(n24876), .B(n24875), .Y(n24878) );
  NOR2XL U11944 ( .A(n24869), .B(n3077), .Y(n24879) );
  NAND2XL U11945 ( .A(n24923), .B(n24922), .Y(n24924) );
  OR2XL U11946 ( .A(n24969), .B(n24968), .Y(n24970) );
  NOR2XL U11947 ( .A(n23369), .B(n23371), .Y(n23382) );
  OAI22XL U11948 ( .A0(n22380), .A1(n22461), .B0(n22265), .B1(n22264), .Y(
        n22464) );
  NOR2XL U11949 ( .A(n22263), .B(n22262), .Y(n22264) );
  NOR2X2 U11950 ( .A(n22389), .B(n22398), .Y(n23272) );
  INVXL U11951 ( .A(n23250), .Y(n23278) );
  INVX1 U11952 ( .A(n23244), .Y(n23346) );
  INVXL U11953 ( .A(n23374), .Y(n23371) );
  NAND2XL U11954 ( .A(n22379), .B(n23337), .Y(n22409) );
  NOR2XL U11955 ( .A(n23329), .B(n22350), .Y(n22379) );
  NAND2XL U11956 ( .A(n23335), .B(n23305), .Y(n22350) );
  OAI22XL U11957 ( .A0(n22462), .A1(n22461), .B0(n22460), .B1(n22459), .Y(
        n23387) );
  NOR2XL U11958 ( .A(n22447), .B(n3082), .Y(n22460) );
  NAND3BXL U11959 ( .AN(n22457), .B(n22456), .C(n3082), .Y(n22458) );
  NAND2XL U11960 ( .A(n21166), .B(target_temp[26]), .Y(n11590) );
  NAND2XL U11961 ( .A(n3111), .B(sigma10[26]), .Y(n11591) );
  NOR2XL U11962 ( .A(n17395), .B(n17399), .Y(n17396) );
  AOI22X2 U11963 ( .A0(n23747), .A1(n3081), .B0(n20690), .B1(n4267), .Y(n24984) );
  INVX1 U11964 ( .A(n24696), .Y(n24188) );
  AOI22XL U11965 ( .A0(n24199), .A1(n4215), .B0(n24179), .B1(n4220), .Y(n24190) );
  AOI22X1 U11966 ( .A0(n23703), .A1(n4267), .B0(n3081), .B1(n5340), .Y(n24224)
         );
  NAND2XL U11967 ( .A(n23784), .B(n25829), .Y(n25703) );
  AND2X1 U11968 ( .A(n23672), .B(n25829), .Y(n25834) );
  AOI22X1 U11969 ( .A0(n20385), .A1(n23833), .B0(n25300), .B1(n23832), .Y(
        n23836) );
  INVXL U11970 ( .A(n23833), .Y(n23830) );
  XOR2XL U11971 ( .A(n25790), .B(n25791), .Y(n25793) );
  NOR2X1 U11972 ( .A(n20783), .B(n20782), .Y(n25722) );
  INVXL U11973 ( .A(n20800), .Y(n20779) );
  AOI22X1 U11974 ( .A0(n20385), .A1(n23805), .B0(n25300), .B1(n23804), .Y(
        n25030) );
  NAND2X1 U11975 ( .A(n23807), .B(n3139), .Y(n5559) );
  NAND2XL U11976 ( .A(n23806), .B(n3455), .Y(n23808) );
  NAND2X1 U11977 ( .A(n20908), .B(n3139), .Y(n5104) );
  INVXL U11978 ( .A(n24091), .Y(n24095) );
  INVX1 U11979 ( .A(n23825), .Y(n23837) );
  NAND2X1 U11980 ( .A(n3455), .B(n20620), .Y(n20621) );
  OAI2BB1X1 U11981 ( .A0N(n23868), .A1N(n23856), .B0(n23855), .Y(n25076) );
  INVXL U11982 ( .A(n25291), .Y(n25287) );
  AND2X2 U11983 ( .A(n20311), .B(n3895), .Y(n4951) );
  OAI2BB1X1 U11984 ( .A0N(n3895), .A1N(n21045), .B0(n13024), .Y(n5968) );
  NAND2X2 U11985 ( .A(n5953), .B(n5952), .Y(n5967) );
  INVX1 U11986 ( .A(n19044), .Y(n4886) );
  INVXL U11987 ( .A(n23515), .Y(n23516) );
  NAND2X1 U11988 ( .A(n5033), .B(n5454), .Y(n5453) );
  NAND2X1 U11989 ( .A(n5450), .B(n5454), .Y(n5449) );
  INVXL U11990 ( .A(n24469), .Y(n24467) );
  INVXL U11991 ( .A(n24502), .Y(n24483) );
  NOR2XL U11992 ( .A(n24586), .B(n24537), .Y(n24539) );
  AOI22XL U11993 ( .A0(n24617), .A1(n24622), .B0(n25290), .B1(n24621), .Y(
        n25521) );
  INVXL U11994 ( .A(n24622), .Y(n24619) );
  INVXL U11995 ( .A(n24658), .Y(n24634) );
  AOI22XL U11996 ( .A0(n24617), .A1(n24703), .B0(n25290), .B1(n24702), .Y(
        n25473) );
  INVXL U11997 ( .A(n24703), .Y(n24700) );
  INVXL U11998 ( .A(n24880), .Y(n21012) );
  XOR2XL U11999 ( .A(n17183), .B(n17406), .Y(n17190) );
  AOI22XL U12000 ( .A0(n22486), .A1(sigma11[25]), .B0(sigma12[25]), .B1(n25754), .Y(n25193) );
  AOI22XL U12001 ( .A0(n22486), .A1(sigma11[29]), .B0(sigma12[29]), .B1(n25754), .Y(n25768) );
  AOI22XL U12002 ( .A0(n25201), .A1(sigma11[24]), .B0(sigma12[24]), .B1(n25754), .Y(n25202) );
  AOI22XL U12003 ( .A0(n22486), .A1(sigma11[3]), .B0(n25754), .B1(sigma12[3]), 
        .Y(n24124) );
  AOI22XL U12004 ( .A0(n22486), .A1(sigma11[17]), .B0(n25754), .B1(sigma12[17]), .Y(n24229) );
  AOI22XL U12005 ( .A0(n22486), .A1(sigma11[22]), .B0(n25754), .B1(sigma12[22]), .Y(n25765) );
  XNOR2XL U12006 ( .A(n25870), .B(n7475), .Y(n7052) );
  INVXL U12007 ( .A(n23158), .Y(n15027) );
  OAI2BB2XL U12008 ( .B0(n22970), .B1(n3225), .A0N(n22987), .A1N(n22969), .Y(
        n22971) );
  XOR2XL U12009 ( .A(n22975), .B(n3055), .Y(n23045) );
  NAND2BXL U12010 ( .AN(n16602), .B(n5847), .Y(n5838) );
  XOR2XL U12011 ( .A(M5_mult_x_15_n1), .B(n16965), .Y(n16575) );
  XNOR2XL U12012 ( .A(n25870), .B(n25881), .Y(n6977) );
  XNOR2XL U12013 ( .A(n25867), .B(n25873), .Y(n7039) );
  XNOR2XL U12014 ( .A(n23221), .B(n25880), .Y(n7026) );
  OAI22XL U12015 ( .A0(n6991), .A1(n25866), .B0(n6990), .B1(n6989), .Y(n7059)
         );
  XNOR2XL U12016 ( .A(n25870), .B(n7569), .Y(n7184) );
  OAI22XL U12017 ( .A0(n9963), .A1(n3182), .B0(n9902), .B1(n3180), .Y(n9897)
         );
  XNOR2XL U12018 ( .A(n9851), .B(n9960), .Y(n9853) );
  XOR2X1 U12019 ( .A(n3108), .B(n4002), .Y(n6137) );
  XNOR2XL U12020 ( .A(n12282), .B(n11499), .Y(n12254) );
  XNOR2X1 U12021 ( .A(n12282), .B(M3_mult_x_15_b_1_), .Y(n12295) );
  NAND2BXL U12022 ( .AN(n3110), .B(n12265), .Y(n12256) );
  XNOR2X1 U12023 ( .A(n12282), .B(n12279), .Y(n12264) );
  INVXL U12024 ( .A(n18235), .Y(n6039) );
  INVXL U12025 ( .A(n6038), .Y(n6036) );
  XOR2XL U12026 ( .A(n5430), .B(M4_U3_U1_or2_inv_0__30_), .Y(n5466) );
  INVXL U12027 ( .A(n8586), .Y(n8333) );
  INVXL U12028 ( .A(n19615), .Y(n19469) );
  INVXL U12029 ( .A(n19676), .Y(n19463) );
  INVXL U12030 ( .A(n15304), .Y(n14999) );
  INVXL U12031 ( .A(n23159), .Y(n15018) );
  INVXL U12032 ( .A(n15283), .Y(n15091) );
  INVXL U12033 ( .A(n15275), .Y(n15088) );
  INVXL U12034 ( .A(n15314), .Y(n15069) );
  AOI22XL U12035 ( .A0(n21507), .A1(n21721), .B0(n21643), .B1(n21697), .Y(
        n21745) );
  INVXL U12036 ( .A(n21683), .Y(n21581) );
  INVXL U12037 ( .A(n21728), .Y(n21534) );
  NAND2XL U12038 ( .A(n21689), .B(n21671), .Y(n21516) );
  NAND2XL U12039 ( .A(n21643), .B(n21458), .Y(n21459) );
  INVXL U12040 ( .A(n21714), .Y(n21458) );
  NAND2XL U12041 ( .A(n21689), .B(n21718), .Y(n21463) );
  INVXL U12042 ( .A(n7165), .Y(n7098) );
  OAI22XL U12043 ( .A0(n7633), .A1(n7061), .B0(n7090), .B1(n7634), .Y(n7096)
         );
  OAI2BB2XL U12044 ( .B0(n22701), .B1(n3225), .A0N(n22987), .A1N(n22700), .Y(
        n22702) );
  XOR2XL U12045 ( .A(n22986), .B(n3056), .Y(n22996) );
  INVXL U12046 ( .A(n22582), .Y(n22583) );
  OAI2BB2XL U12047 ( .B0(n22709), .B1(n3225), .A0N(n22987), .A1N(n22708), .Y(
        n22710) );
  XOR2XL U12048 ( .A(n22714), .B(n22713), .Y(n22722) );
  NAND2XL U12049 ( .A(n22892), .B(n22987), .Y(n4708) );
  OAI22X1 U12050 ( .A0(n7511), .A1(n6433), .B0(n7512), .B1(n6379), .Y(n6407)
         );
  XNOR2XL U12051 ( .A(M0_b_1_), .B(n25869), .Y(n6410) );
  NOR2BXL U12052 ( .AN(n6944), .B(n6990), .Y(n6566) );
  NAND2XL U12053 ( .A(n6845), .B(M0_b_1_), .Y(n6565) );
  NAND2BXL U12054 ( .AN(n6944), .B(n21054), .Y(n6563) );
  NAND2BXL U12055 ( .AN(n6944), .B(n3209), .Y(n6549) );
  CMPR32X1 U12056 ( .A(n6619), .B(n6618), .C(n6617), .CO(n6624), .S(n6626) );
  NOR2BXL U12057 ( .AN(n6944), .B(n6608), .Y(n6619) );
  INVXL U12058 ( .A(n6499), .Y(n5632) );
  OAI21XL U12059 ( .A0(n7093), .A1(n6500), .B0(n5635), .Y(n5634) );
  NAND2BXL U12060 ( .AN(n6474), .B(n6293), .Y(n5635) );
  OAI22XL U12061 ( .A0(n6845), .A1(n6362), .B0(n6321), .B1(n6843), .Y(n6329)
         );
  OAI22XL U12062 ( .A0(n6613), .A1(n6393), .B0(n6608), .B1(n6322), .Y(n6328)
         );
  CMPR32X1 U12063 ( .A(n7113), .B(n7112), .C(n7111), .CO(n7141), .S(n7108) );
  OAI22XL U12064 ( .A0(n7511), .A1(n7050), .B0(n7512), .B1(n7091), .Y(n7112)
         );
  NAND2BXL U12065 ( .AN(n16630), .B(n3044), .Y(n5836) );
  NAND2BXL U12066 ( .AN(n3110), .B(n3047), .Y(n16630) );
  OAI22XL U12067 ( .A0(n16640), .A1(n5835), .B0(n16629), .B1(n16704), .Y(
        n16641) );
  OAI22XL U12068 ( .A0(n16638), .A1(n16628), .B0(n16637), .B1(n16475), .Y(
        n16642) );
  NAND2BXL U12069 ( .AN(n16703), .B(n5847), .Y(n5843) );
  XNOR2XL U12070 ( .A(n16614), .B(n11499), .Y(n16569) );
  XNOR2XL U12071 ( .A(n16614), .B(n16884), .Y(n16473) );
  OAI22XL U12072 ( .A0(n7093), .A1(n7027), .B0(n7094), .B1(n3209), .Y(n7046)
         );
  XNOR2XL U12073 ( .A(n25867), .B(n25874), .Y(n6978) );
  XNOR2XL U12074 ( .A(M0_b_9_), .B(n23221), .Y(n6988) );
  XNOR2XL U12075 ( .A(n25869), .B(n7569), .Y(n7028) );
  XNOR2XL U12076 ( .A(n25867), .B(n25872), .Y(n7088) );
  NAND2BXL U12077 ( .AN(n7089), .B(n3188), .Y(n5116) );
  XNOR2XL U12078 ( .A(n25870), .B(n25879), .Y(n7148) );
  XNOR2XL U12079 ( .A(n25870), .B(n7621), .Y(n7292) );
  XNOR2XL U12080 ( .A(n25869), .B(n25874), .Y(n7466) );
  XNOR2X1 U12081 ( .A(n25869), .B(n7646), .Y(n7222) );
  XNOR2XL U12082 ( .A(n25869), .B(n25876), .Y(n7185) );
  XNOR2X1 U12083 ( .A(M2_mult_x_15_n43), .B(n10386), .Y(n9361) );
  NAND2XL U12084 ( .A(n9966), .B(n10159), .Y(n6059) );
  XNOR2X1 U12085 ( .A(M2_a_17_), .B(n10514), .Y(n10301) );
  XNOR2XL U12086 ( .A(n9904), .B(n9874), .Y(n9873) );
  ADDHXL U12087 ( .A(n9917), .B(n9916), .CO(n9918), .S(n9910) );
  OAI22XL U12088 ( .A0(n9963), .A1(n9902), .B0(n9913), .B1(n3180), .Y(n9917)
         );
  OAI22XL U12089 ( .A0(n9983), .A1(n9903), .B0(n9981), .B1(n9915), .Y(n9916)
         );
  XNOR2XL U12090 ( .A(n9904), .B(n9960), .Y(n9903) );
  XNOR2XL U12091 ( .A(n9841), .B(n9960), .Y(n9834) );
  XNOR2X1 U12092 ( .A(n9904), .B(n9836), .Y(n9840) );
  XNOR2X1 U12093 ( .A(M2_mult_x_15_a_1_), .B(n10514), .Y(n9631) );
  NOR2XL U12094 ( .A(n9222), .B(n3180), .Y(n9224) );
  OAI22X1 U12095 ( .A0(n10660), .A1(n3182), .B0(n3178), .B1(n9892), .Y(n9225)
         );
  NOR2BXL U12096 ( .AN(n3110), .B(n12222), .Y(n12259) );
  XNOR2XL U12097 ( .A(n12519), .B(n11499), .Y(n12066) );
  OAI22X1 U12098 ( .A0(n12340), .A1(n4877), .B0(n12338), .B1(n12064), .Y(
        n12097) );
  NOR2BXL U12099 ( .AN(n3110), .B(n12718), .Y(n12098) );
  OAI22XL U12100 ( .A0(n12597), .A1(n12072), .B0(n12595), .B1(n12009), .Y(
        n12069) );
  NAND2BXL U12101 ( .AN(n3110), .B(M3_mult_x_15_a_17_), .Y(n12032) );
  XNOR2XL U12102 ( .A(n12282), .B(n3198), .Y(n12010) );
  XNOR2X1 U12103 ( .A(n12594), .B(n3197), .Y(n12009) );
  XOR2XL U12104 ( .A(n5430), .B(n12522), .Y(n5516) );
  XNOR2XL U12105 ( .A(n25884), .B(n11499), .Y(n12027) );
  XNOR2XL U12106 ( .A(n13864), .B(n4807), .Y(n13053) );
  XNOR2XL U12107 ( .A(n13919), .B(n13693), .Y(n13065) );
  ADDHXL U12108 ( .A(n13118), .B(n13117), .CO(n13119), .S(n13111) );
  OAI22XL U12109 ( .A0(n13790), .A1(n13720), .B0(n13106), .B1(n13721), .Y(
        n13118) );
  OAI22XL U12110 ( .A0(n13114), .A1(n3181), .B0(n13107), .B1(n13532), .Y(
        n13117) );
  NAND2BXL U12111 ( .AN(n13049), .B(n25860), .Y(n13106) );
  NOR2BXL U12112 ( .AN(n13049), .B(n13972), .Y(n13088) );
  OAI22XL U12113 ( .A0(n13085), .A1(n13790), .B0(n13074), .B1(n13721), .Y(
        n13087) );
  OAI22XL U12114 ( .A0(n13056), .A1(n3181), .B0(n13075), .B1(n13532), .Y(
        n13072) );
  NAND2BXL U12115 ( .AN(n13049), .B(n4807), .Y(n13050) );
  XNOR2XL U12116 ( .A(n13919), .B(n13844), .Y(n13156) );
  XNOR2XL U12117 ( .A(n14027), .B(n13844), .Y(n13206) );
  XNOR2XL U12118 ( .A(n14028), .B(n13844), .Y(n13168) );
  XNOR2XL U12119 ( .A(n4567), .B(n25860), .Y(n13208) );
  XNOR2XL U12120 ( .A(n4565), .B(n13844), .Y(n13220) );
  XOR2XL U12121 ( .A(n13769), .B(n5512), .Y(n13259) );
  XNOR2XL U12122 ( .A(n13049), .B(n25862), .Y(n13262) );
  XNOR2XL U12123 ( .A(n4567), .B(n13844), .Y(n13267) );
  NAND2BXL U12124 ( .AN(n13049), .B(n25862), .Y(n13281) );
  XNOR2XL U12125 ( .A(n14117), .B(n4848), .Y(n13314) );
  XOR2XL U12126 ( .A(n13863), .B(n5512), .Y(n13317) );
  XNOR2XL U12127 ( .A(n13919), .B(M1_b_11_), .Y(n13318) );
  NAND2X1 U12128 ( .A(n3123), .B(w1[133]), .Y(n5262) );
  NAND2X1 U12129 ( .A(target_temp[12]), .B(n9164), .Y(n5491) );
  OAI21XL U12130 ( .A0(n25243), .A1(n26232), .B0(n11516), .Y(M1_a_9_) );
  XNOR2X1 U12131 ( .A(n18006), .B(n3201), .Y(n17904) );
  XNOR2XL U12132 ( .A(n18604), .B(n2978), .Y(n17900) );
  XNOR2X1 U12133 ( .A(n18604), .B(M3_mult_x_15_b_1_), .Y(n17899) );
  XNOR2XL U12134 ( .A(n3206), .B(n11499), .Y(n18138) );
  XNOR2XL U12135 ( .A(n18006), .B(n11499), .Y(n18175) );
  XNOR2X1 U12136 ( .A(n18006), .B(M3_mult_x_15_b_3_), .Y(n18176) );
  XNOR2XL U12137 ( .A(n3206), .B(n12271), .Y(n18178) );
  XOR2XL U12138 ( .A(M3_mult_x_15_b_1_), .B(n18169), .Y(n18179) );
  OAI22XL U12139 ( .A0(n18242), .A1(n18169), .B0(n18168), .B1(n18167), .Y(
        n18171) );
  NOR2BXL U12140 ( .AN(n2978), .B(n18168), .Y(n18160) );
  OAI22XL U12141 ( .A0(n18177), .A1(n2978), .B0(M3_mult_x_15_b_1_), .B1(n18223), .Y(n18159) );
  NAND2BXL U12142 ( .AN(n2978), .B(n18006), .Y(n18157) );
  ADDHXL U12143 ( .A(n18181), .B(n18180), .CO(n18182), .S(n18172) );
  OAI22XL U12144 ( .A0(n18242), .A1(n18166), .B0(n18168), .B1(n18179), .Y(
        n18180) );
  OAI22XL U12145 ( .A0(n18177), .A1(n18165), .B0(n18176), .B1(n18223), .Y(
        n18181) );
  XNOR2XL U12146 ( .A(n3206), .B(n2978), .Y(n18166) );
  CMPR32X1 U12147 ( .A(n18145), .B(n18144), .C(n18143), .CO(n18136), .S(n18146) );
  XOR2X1 U12148 ( .A(n18142), .B(n2974), .Y(n5918) );
  XOR2X1 U12149 ( .A(M3_mult_x_15_n1682), .B(n3189), .Y(n5820) );
  XNOR2XL U12150 ( .A(n18468), .B(n2978), .Y(n17969) );
  OR2X2 U12151 ( .A(n17975), .B(n18235), .Y(n5459) );
  XNOR2XL U12152 ( .A(n18006), .B(n18611), .Y(n17994) );
  XNOR2XL U12153 ( .A(n14235), .B(n4848), .Y(n13477) );
  NOR2XL U12154 ( .A(n3214), .B(n3181), .Y(n13691) );
  OAI22XL U12155 ( .A0(n13694), .A1(n13790), .B0(n13721), .B1(n13693), .Y(
        n13715) );
  OAI22XL U12156 ( .A0(n2993), .A1(n13864), .B0(n14356), .B1(n13863), .Y(
        n13716) );
  INVXL U12157 ( .A(n13864), .Y(n13768) );
  OAI22XL U12158 ( .A0(n2993), .A1(n25865), .B0(n14356), .B1(n13919), .Y(
        n13862) );
  XNOR2XL U12159 ( .A(n14195), .B(n25862), .Y(n13838) );
  OAI21XL U12160 ( .A0(n3092), .A1(n8532), .B0(n8301), .Y(n8363) );
  INVXL U12161 ( .A(n8554), .Y(n8336) );
  INVXL U12162 ( .A(n23179), .Y(n8281) );
  AOI2BB2XL U12163 ( .B0(n8371), .B1(n3157), .A0N(n3157), .A1N(n8433), .Y(
        n8512) );
  INVXL U12164 ( .A(n19643), .Y(n19466) );
  NAND2XL U12165 ( .A(n19564), .B(n19386), .Y(n19387) );
  INVXL U12166 ( .A(n15118), .Y(n14992) );
  NAND2XL U12167 ( .A(n21643), .B(n21471), .Y(n21472) );
  INVXL U12168 ( .A(n21699), .Y(n21471) );
  AOI22XL U12169 ( .A0(n3095), .A1(n21661), .B0(n21629), .B1(n21580), .Y(
        n21798) );
  INVXL U12170 ( .A(n15176), .Y(n15223) );
  INVXL U12171 ( .A(n15171), .Y(n15192) );
  INVXL U12172 ( .A(n15105), .Y(n15151) );
  NAND2XL U12173 ( .A(n3038), .B(n15279), .Y(n15081) );
  INVXL U12174 ( .A(n15288), .Y(n15139) );
  NAND2XL U12175 ( .A(n21580), .B(n21540), .Y(n21541) );
  INVXL U12176 ( .A(n21588), .Y(n21540) );
  NAND2XL U12177 ( .A(n21580), .B(n21564), .Y(n21565) );
  AOI22XL U12178 ( .A0(n3095), .A1(n21591), .B0(n21590), .B1(n21580), .Y(
        n21781) );
  INVXL U12179 ( .A(n21589), .Y(n21590) );
  NAND2XL U12180 ( .A(n21580), .B(n21592), .Y(n21593) );
  NAND2XL U12181 ( .A(n21580), .B(n21586), .Y(n21587) );
  INVXL U12182 ( .A(n21585), .Y(n21586) );
  NAND2XL U12183 ( .A(n21580), .B(n21547), .Y(n21548) );
  INVXL U12184 ( .A(n21594), .Y(n21547) );
  NAND2XL U12185 ( .A(n21741), .B(n3171), .Y(n21595) );
  AOI2BB2XL U12186 ( .B0(n21855), .B1(n3096), .A0N(n3096), .A1N(n21795), .Y(
        n21618) );
  XNOR2XL U12187 ( .A(n23221), .B(n25874), .Y(n7536) );
  XNOR2XL U12188 ( .A(n23221), .B(n25873), .Y(n7547) );
  XNOR2XL U12189 ( .A(n25870), .B(n25875), .Y(n7546) );
  INVXL U12190 ( .A(n22928), .Y(n22701) );
  XNOR2XL U12191 ( .A(n23221), .B(n7800), .Y(n7570) );
  XNOR2XL U12192 ( .A(n23221), .B(n25872), .Y(n7589) );
  XNOR2XL U12193 ( .A(n25870), .B(n25874), .Y(n7563) );
  XNOR2XL U12194 ( .A(n25870), .B(n25873), .Y(n7588) );
  INVXL U12195 ( .A(n22988), .Y(n22981) );
  XNOR2XL U12196 ( .A(n25869), .B(n25872), .Y(n7555) );
  XNOR2XL U12197 ( .A(n25869), .B(n7800), .Y(n7531) );
  XNOR2XL U12198 ( .A(n25870), .B(n7646), .Y(n7532) );
  XNOR2X1 U12199 ( .A(n23221), .B(n7646), .Y(n7459) );
  XOR2XL U12200 ( .A(n22699), .B(n3058), .Y(n22726) );
  AOI222XL U12201 ( .A0(n22928), .A1(n10749), .B0(n22700), .B1(n3116), .C0(
        n22927), .C1(n22987), .Y(n22697) );
  AOI222XL U12202 ( .A0(n22953), .A1(n11074), .B0(n10797), .B1(n3219), .C0(
        n22952), .C1(n11073), .Y(n22799) );
  NOR2XL U12203 ( .A(n10769), .B(n23002), .Y(n10812) );
  NAND2XL U12204 ( .A(n23002), .B(n10749), .Y(n10822) );
  NAND2XL U12205 ( .A(n10769), .B(n23002), .Y(n10813) );
  OAI22XL U12206 ( .A0(n23193), .A1(n26225), .B0(n9107), .B1(n25942), .Y(
        n11144) );
  OAI22XL U12207 ( .A0(n23193), .A1(n26228), .B0(n9107), .B1(n25941), .Y(
        n11146) );
  INVXL U12208 ( .A(n5576), .Y(M0_U4_U1_enc_tree_1__1__28_) );
  NOR2XL U12209 ( .A(M0_a_7_), .B(M0_a_6_), .Y(M0_U3_U1_enc_tree_1__1__24_) );
  NOR2XL U12210 ( .A(n5398), .B(M0_a_15_), .Y(M0_U3_U1_enc_tree_1__1__16_) );
  OAI22XL U12211 ( .A0(n7287), .A1(n6397), .B0(n6364), .B1(n7288), .Y(n6405)
         );
  NOR2BXL U12212 ( .AN(n6944), .B(n7094), .Y(n6581) );
  OAI22XL U12213 ( .A0(n6571), .A1(n6991), .B0(n6561), .B1(n6602), .Y(n6579)
         );
  OAI22XL U12214 ( .A0(n6572), .A1(n6845), .B0(n6560), .B1(n6843), .Y(n6580)
         );
  NAND2BXL U12215 ( .AN(n6944), .B(n25866), .Y(n6569) );
  XNOR2XL U12216 ( .A(n25867), .B(n6944), .Y(n6607) );
  ADDFX2 U12217 ( .A(n6599), .B(n6600), .CI(n6598), .CO(n6649), .S(n6657) );
  NOR2BXL U12218 ( .AN(n6944), .B(n7288), .Y(n6600) );
  ADDFX2 U12219 ( .A(n6648), .B(n6647), .CI(n6646), .CO(n6653), .S(n6655) );
  OAI22XL U12220 ( .A0(n6614), .A1(n6613), .B0(n6612), .B1(n7146), .Y(n6646)
         );
  CMPR32X1 U12221 ( .A(n6512), .B(n6511), .C(n6510), .CO(n6504), .S(n6642) );
  OAI22XL U12222 ( .A0(n6503), .A1(n7287), .B0(n6493), .B1(n7288), .Y(n6511)
         );
  CMPR32X1 U12223 ( .A(n6458), .B(n6457), .C(n6456), .CO(n6453), .S(n6678) );
  NOR2BXL U12224 ( .AN(n6944), .B(n3046), .Y(n6458) );
  NAND2BXL U12225 ( .AN(n6944), .B(n25870), .Y(n6315) );
  XNOR2XL U12226 ( .A(n25870), .B(n6944), .Y(n6345) );
  CLKINVX3 U12227 ( .A(n5583), .Y(n6608) );
  AOI22XL U12228 ( .A0(n7389), .A1(target_temp[10]), .B0(in_valid_d), .B1(
        w1[10]), .Y(n6228) );
  AOI22X1 U12229 ( .A0(n7389), .A1(target_temp[17]), .B0(n3123), .B1(w1[17]), 
        .Y(n6237) );
  OAI21XL U12230 ( .A0(n6274), .A1(n26224), .B0(n6253), .Y(M0_b_15_) );
  AOI21XL U12231 ( .A0(n6733), .A1(y10[1]), .B0(n25139), .Y(n6278) );
  NOR2BXL U12232 ( .AN(n5983), .B(M3_a_9_), .Y(M3_U3_U1_enc_tree_1__1__22_) );
  INVXL U12233 ( .A(M3_U3_U1_enc_tree_1__1__28_), .Y(M3_U3_U1_or2_inv_1__28_)
         );
  INVXL U12234 ( .A(M3_U3_U1_or2_tree_1__2__24_), .Y(M3_U3_U1_or2_inv_1__24_)
         );
  NOR2XL U12235 ( .A(M3_mult_x_15_n61), .B(M3_a_20_), .Y(
        M3_U3_U1_enc_tree_1__1__10_) );
  INVXL U12236 ( .A(M3_U3_U1_enc_tree_2__2__24_), .Y(M3_U3_U1_or2_inv_2__24_)
         );
  NOR2XL U12237 ( .A(M3_mult_x_15_a_17_), .B(M3_a_16_), .Y(
        M3_U3_U1_enc_tree_1__1__14_) );
  ADDFX2 U12238 ( .A(n16612), .B(n16610), .CI(n16611), .CO(n16661), .S(n16660)
         );
  NAND2BXL U12239 ( .AN(n16613), .B(n5847), .Y(n5840) );
  NOR2BXL U12240 ( .AN(n3110), .B(n16699), .Y(n16653) );
  OAI22XL U12241 ( .A0(n16701), .A1(n16616), .B0(n16699), .B1(n16615), .Y(
        n16649) );
  XNOR2XL U12242 ( .A(n16614), .B(n3110), .Y(n16616) );
  NAND2BXL U12243 ( .AN(n16573), .B(n5847), .Y(n5841) );
  OAI21X1 U12244 ( .A0(n16532), .A1(n5835), .B0(n5842), .Y(n16544) );
  OAI22XL U12245 ( .A0(n16701), .A1(n16698), .B0(n16699), .B1(n6145), .Y(
        n16681) );
  OAI21XL U12246 ( .A0(n16687), .A1(n16942), .B0(n5733), .Y(n16680) );
  CMPR32X1 U12247 ( .A(n16707), .B(n16706), .C(n16705), .CO(n16744), .S(n16739) );
  ADDFX2 U12248 ( .A(n16738), .B(n16736), .CI(n16737), .CO(n16546), .S(n16747)
         );
  OAI21XL U12249 ( .A0(n16516), .A1(n16688), .B0(n5731), .Y(n16738) );
  NOR2X1 U12250 ( .A(n5548), .B(n5547), .Y(n5546) );
  NOR2XL U12251 ( .A(n16401), .B(n16942), .Y(n5547) );
  NOR2XL U12252 ( .A(n16353), .B(n16688), .Y(n5548) );
  CMPR32X1 U12253 ( .A(n16489), .B(n16488), .C(n16487), .CO(n16486), .S(n16557) );
  XNOR2XL U12254 ( .A(n3211), .B(M3_mult_x_15_b_2_), .Y(n16348) );
  XOR2XL U12255 ( .A(n17039), .B(n5705), .Y(n5704) );
  OAI21X1 U12256 ( .A0(n5835), .A1(n16344), .B0(n5860), .Y(n5859) );
  OAI22X1 U12257 ( .A0(n16701), .A1(n16361), .B0(n16699), .B1(n16360), .Y(
        n16371) );
  OAI22XL U12258 ( .A0(n16942), .A1(n16359), .B0(n16688), .B1(n16379), .Y(
        n16372) );
  XOR2XL U12259 ( .A(n6124), .B(n17039), .Y(n5706) );
  XNOR2XL U12260 ( .A(n16614), .B(n12701), .Y(n16360) );
  XNOR2XL U12261 ( .A(n16614), .B(n3198), .Y(n16328) );
  XOR2X1 U12262 ( .A(n12279), .B(n3212), .Y(n5693) );
  XNOR2XL U12263 ( .A(n3211), .B(M3_mult_x_15_b_6_), .Y(n16103) );
  OAI22XL U12264 ( .A0(n16942), .A1(n16379), .B0(n16688), .B1(n16378), .Y(
        n16440) );
  OAI22X2 U12265 ( .A0(n17060), .A1(n16377), .B0(n17061), .B1(n5706), .Y(
        n16427) );
  OAI22X2 U12266 ( .A0(n17074), .A1(n16376), .B0(n16375), .B1(n16374), .Y(
        n16428) );
  XNOR2X1 U12267 ( .A(n5677), .B(n3110), .Y(n16376) );
  NOR2X1 U12268 ( .A(n16373), .B(n16939), .Y(n5806) );
  NOR2BXL U12269 ( .AN(n3110), .B(n16317), .Y(n16426) );
  NOR2XL U12270 ( .A(n3203), .B(M5_a_10_), .Y(M5_U3_U1_enc_tree_1__1__20_) );
  INVXL U12271 ( .A(M5_U3_U1_enc_tree_1__1__28_), .Y(M5_U3_U1_or2_inv_1__28_)
         );
  INVXL U12272 ( .A(M5_U3_U1_or2_tree_1__2__24_), .Y(M5_U3_U1_or2_inv_1__24_)
         );
  INVXL U12273 ( .A(M5_U3_U1_enc_tree_2__2__24_), .Y(M5_U3_U1_or2_inv_2__24_)
         );
  NAND2XL U12274 ( .A(n11188), .B(n11187), .Y(n21063) );
  NAND2XL U12275 ( .A(w2[77]), .B(valid[0]), .Y(n11187) );
  NAND2XL U12276 ( .A(w2[45]), .B(n23973), .Y(n11188) );
  NAND2XL U12277 ( .A(n11190), .B(n11189), .Y(n21062) );
  NAND2XL U12278 ( .A(w2[76]), .B(valid[0]), .Y(n11189) );
  NAND2XL U12279 ( .A(w2[44]), .B(n23973), .Y(n11190) );
  NAND2XL U12280 ( .A(n11180), .B(n11179), .Y(n21059) );
  NAND2XL U12281 ( .A(w2[80]), .B(valid[0]), .Y(n11179) );
  NAND2XL U12282 ( .A(w2[48]), .B(n3501), .Y(n11180) );
  NAND2XL U12283 ( .A(w2[78]), .B(valid[0]), .Y(n11184) );
  NAND2XL U12284 ( .A(w2[46]), .B(n23973), .Y(n11185) );
  NAND2XL U12285 ( .A(n11183), .B(n11182), .Y(n21058) );
  NAND2XL U12286 ( .A(w2[79]), .B(valid[0]), .Y(n11182) );
  NAND2XL U12287 ( .A(w2[47]), .B(n23973), .Y(n11183) );
  OAI22XL U12288 ( .A0(n11057), .A1(n26214), .B0(n9107), .B1(n25948), .Y(
        n11152) );
  OAI22XL U12289 ( .A0(n11057), .A1(n26215), .B0(n9107), .B1(n25947), .Y(
        n11154) );
  XNOR2X1 U12290 ( .A(n17039), .B(n16965), .Y(n5642) );
  XNOR2X1 U12291 ( .A(n3203), .B(n3196), .Y(n16200) );
  NAND2XL U12292 ( .A(n8482), .B(n8313), .Y(n8314) );
  INVXL U12293 ( .A(n8407), .Y(n8421) );
  INVXL U12294 ( .A(n8424), .Y(n8460) );
  NAND2XL U12295 ( .A(n7077), .B(n7076), .Y(n7127) );
  NAND2XL U12296 ( .A(n7075), .B(n7074), .Y(n7076) );
  XNOR2XL U12297 ( .A(n25867), .B(n25875), .Y(n6931) );
  CMPR32X1 U12298 ( .A(n7144), .B(n7143), .C(n7142), .CO(n7200), .S(n7154) );
  ADDFX2 U12299 ( .A(n7300), .B(n7299), .CI(n7298), .CO(n7476), .S(n7302) );
  XNOR2XL U12300 ( .A(n25870), .B(n25878), .Y(n7227) );
  OAI22X1 U12301 ( .A0(n10660), .A1(n10311), .B0(n3178), .B1(n10342), .Y(n5543) );
  INVXL U12302 ( .A(n10312), .Y(n10171) );
  OAI22XL U12303 ( .A0(n10532), .A1(n9216), .B0(n9215), .B1(n9362), .Y(n9354)
         );
  INVXL U12304 ( .A(n9478), .Y(n5301) );
  INVXL U12305 ( .A(n9836), .Y(n9359) );
  XNOR2X1 U12306 ( .A(n10494), .B(n10386), .Y(n9581) );
  XNOR2XL U12307 ( .A(n10337), .B(n5298), .Y(n10330) );
  OAI22XL U12308 ( .A0(n4570), .A1(n9700), .B0(n10403), .B1(n9666), .Y(n9696)
         );
  NOR2BX1 U12309 ( .AN(n9960), .B(n10496), .Y(n9698) );
  OAI22XL U12310 ( .A0(n9983), .A1(n9914), .B0(n9981), .B1(n9885), .Y(n9925)
         );
  OAI22XL U12311 ( .A0(n9979), .A1(n9888), .B0(n9977), .B1(n9887), .Y(n9924)
         );
  XNOR2XL U12312 ( .A(n9886), .B(n9960), .Y(n9888) );
  OAI22XL U12313 ( .A0(n9983), .A1(n9915), .B0(n9981), .B1(n9914), .Y(n9926)
         );
  OAI22XL U12314 ( .A0(n9963), .A1(n9913), .B0(n9912), .B1(n3180), .Y(n9927)
         );
  OAI22XL U12315 ( .A0(n9979), .A1(n9721), .B0(n9977), .B1(n9673), .Y(n9714)
         );
  OAI22X1 U12316 ( .A0(n9983), .A1(n9706), .B0(n9981), .B1(n9668), .Y(n9710)
         );
  OAI22XL U12317 ( .A0(n9966), .A1(n9699), .B0(n10159), .B1(n9667), .Y(n9711)
         );
  INVXL U12318 ( .A(n5188), .Y(n5186) );
  OAI22X1 U12319 ( .A0(n9966), .A1(n9798), .B0(n10159), .B1(n9753), .Y(n9797)
         );
  OAI22X1 U12320 ( .A0(n9983), .A1(n9668), .B0(n9981), .B1(n9640), .Y(n9671)
         );
  XNOR2X1 U12321 ( .A(n25885), .B(n3182), .Y(n9396) );
  NOR2XL U12322 ( .A(n10337), .B(M2_b_15_), .Y(M2_U4_U1_enc_tree_1__1__16_) );
  NOR2XL U12323 ( .A(n10341), .B(n10342), .Y(M2_U4_U1_enc_tree_1__1__20_) );
  NOR2XL U12324 ( .A(M2_a_8_), .B(n9841), .Y(M2_U3_U1_enc_tree_1__1__22_) );
  CMPR32X1 U12325 ( .A(n9275), .B(n9274), .C(n9273), .CO(n9351), .S(n9271) );
  INVXL U12326 ( .A(n10341), .Y(n5377) );
  XNOR2X1 U12327 ( .A(M2_a_8_), .B(n9843), .Y(n9214) );
  OAI22XL U12328 ( .A0(n9551), .A1(n9227), .B0(n9838), .B1(n9207), .Y(n9244)
         );
  OAI22X1 U12329 ( .A0(n10517), .A1(n9240), .B0(n10533), .B1(n9204), .Y(n9243)
         );
  XNOR2XL U12330 ( .A(n12758), .B(n11499), .Y(n11690) );
  OAI22XL U12331 ( .A0(n12352), .A1(n12172), .B0(n12222), .B1(n12162), .Y(
        n12183) );
  OAI22XL U12332 ( .A0(n12635), .A1(n12164), .B0(n12513), .B1(n12163), .Y(
        n12182) );
  OAI22XL U12333 ( .A0(n12352), .A1(n12162), .B0(n12222), .B1(n12131), .Y(
        n12167) );
  CMPR32X1 U12334 ( .A(n12199), .B(n12198), .C(n12197), .CO(n12191), .S(n12387) );
  NAND2BXL U12335 ( .AN(n3110), .B(n25884), .Y(n12095) );
  OAI22XL U12336 ( .A0(n12340), .A1(n12120), .B0(n12338), .B1(n4877), .Y(
        n12118) );
  XNOR2X1 U12337 ( .A(n12519), .B(n5430), .Y(n11852) );
  NAND2BXL U12338 ( .AN(n3110), .B(n12732), .Y(n11849) );
  XNOR2X1 U12339 ( .A(n12732), .B(M3_mult_x_15_b_1_), .Y(n12002) );
  XNOR2XL U12340 ( .A(n14288), .B(n25862), .Y(n14075) );
  XNOR2XL U12341 ( .A(n14306), .B(n14156), .Y(n14070) );
  XNOR2XL U12342 ( .A(n14156), .B(n14357), .Y(n5510) );
  XNOR2X1 U12343 ( .A(n14307), .B(n25862), .Y(n14089) );
  XNOR2X1 U12344 ( .A(n18604), .B(n3201), .Y(n18499) );
  XNOR2X1 U12345 ( .A(n18150), .B(M3_mult_x_15_b_12_), .Y(n17941) );
  XNOR2X1 U12346 ( .A(M3_mult_x_15_b_13_), .B(n18150), .Y(n5815) );
  XNOR2X1 U12347 ( .A(n18500), .B(n3197), .Y(n17879) );
  XNOR2XL U12348 ( .A(n18638), .B(n2978), .Y(n17873) );
  XNOR2X1 U12349 ( .A(n18638), .B(M3_mult_x_15_b_1_), .Y(n17871) );
  NOR2BXL U12350 ( .AN(n13049), .B(n13843), .Y(n13129) );
  OAI22XL U12351 ( .A0(n13116), .A1(n13790), .B0(n13115), .B1(n13721), .Y(
        n13127) );
  OAI22XL U12352 ( .A0(n13094), .A1(n13899), .B0(n13093), .B1(n2997), .Y(
        n13125) );
  INVXL U12353 ( .A(n5164), .Y(n5162) );
  CMPR32X1 U12354 ( .A(n13395), .B(n13394), .C(n13393), .CO(n13454), .S(n13405) );
  OAI22XL U12355 ( .A0(n13401), .A1(n14120), .B0(n13359), .B1(n14121), .Y(
        n13393) );
  NAND2X1 U12356 ( .A(in_valid_d), .B(w1[137]), .Y(n5166) );
  XNOR2XL U12357 ( .A(n14117), .B(n14030), .Y(n13481) );
  XNOR2XL U12358 ( .A(n13919), .B(n25862), .Y(n13483) );
  OAI22XL U12359 ( .A0(n14267), .A1(n14282), .B0(n13429), .B1(n14251), .Y(
        n13499) );
  OAI22XL U12360 ( .A0(n13476), .A1(n3181), .B0(n13430), .B1(n13532), .Y(
        n13498) );
  NAND2BXL U12361 ( .AN(n13049), .B(n25863), .Y(n13429) );
  XOR2XL U12362 ( .A(n14028), .B(n5512), .Y(n13449) );
  XNOR2X1 U12363 ( .A(n14265), .B(n13693), .Y(n13482) );
  XNOR2XL U12364 ( .A(n14266), .B(n13693), .Y(n13450) );
  NOR2XL U12365 ( .A(n4807), .B(M1_b_6_), .Y(M1_U4_U1_enc_tree_1__1__24_) );
  NOR2XL U12366 ( .A(n13693), .B(M1_b_2_), .Y(M1_U4_U1_enc_tree_1__1__28_) );
  INVXL U12367 ( .A(M1_U4_U1_enc_tree_2__2__24_), .Y(M1_U4_U1_or2_inv_2__24_)
         );
  INVXL U12368 ( .A(M1_U3_U1_enc_tree_2__2__24_), .Y(M1_U3_U1_or2_inv_2__24_)
         );
  XNOR2XL U12369 ( .A(n14196), .B(n25863), .Y(n13973) );
  XNOR2XL U12370 ( .A(n14117), .B(n25863), .Y(n13917) );
  INVXL U12371 ( .A(n14028), .Y(n13969) );
  CMPR32X1 U12372 ( .A(n14050), .B(n14049), .C(n14048), .CO(n14106), .S(n14042) );
  OAI22XL U12373 ( .A0(n14025), .A1(n14282), .B0(n14059), .B1(n14251), .Y(
        n14048) );
  XNOR2XL U12374 ( .A(n14306), .B(n25862), .Y(n14134) );
  XNOR2XL U12375 ( .A(n5677), .B(n11499), .Y(n16007) );
  OAI22XL U12376 ( .A0(n18239), .A1(n18120), .B0(n18238), .B1(n18104), .Y(
        n18122) );
  OAI22XL U12377 ( .A0(n18242), .A1(n18108), .B0(n18168), .B1(n18241), .Y(
        n18251) );
  OAI22XL U12378 ( .A0(n18239), .A1(n18005), .B0(n18238), .B1(n17992), .Y(
        n18022) );
  OAI21XL U12379 ( .A0(n18235), .A1(n5460), .B0(n5457), .Y(n18045) );
  OAI22XL U12380 ( .A0(n18177), .A1(n18067), .B0(n18049), .B1(n18223), .Y(
        n18070) );
  NOR2BXL U12381 ( .AN(n2978), .B(n5893), .Y(n18071) );
  OAI22X1 U12382 ( .A0(n18083), .A1(n6026), .B0(n18429), .B1(n18050), .Y(
        n18069) );
  XOR2X1 U12383 ( .A(n2974), .B(n18603), .Y(n17693) );
  NAND2X1 U12384 ( .A(n11538), .B(n11537), .Y(M1_b_18_) );
  NAND2X1 U12385 ( .A(n3123), .B(w1[144]), .Y(n11534) );
  XNOR2XL U12386 ( .A(n14307), .B(n25863), .Y(n14210) );
  XNOR2XL U12387 ( .A(n14306), .B(n14228), .Y(n14190) );
  XOR2XL U12388 ( .A(n14196), .B(n6210), .Y(n13540) );
  OAI21X1 U12389 ( .A0(n14157), .A1(n13728), .B0(n5503), .Y(n13795) );
  OAI22XL U12390 ( .A0(n13729), .A1(n14044), .B0(n13779), .B1(n13974), .Y(
        n13794) );
  INVXL U12391 ( .A(n8614), .Y(n8493) );
  INVXL U12392 ( .A(n19648), .Y(n19460) );
  INVXL U12393 ( .A(n19659), .Y(n19458) );
  NAND2XL U12394 ( .A(n20374), .B(n8275), .Y(n8276) );
  AOI2BB2XL U12395 ( .B0(n3040), .B1(n8478), .A0N(n8482), .A1N(n8497), .Y(
        n8572) );
  INVXL U12396 ( .A(n8540), .Y(n8393) );
  INVXL U12397 ( .A(n8536), .Y(n8391) );
  INVXL U12398 ( .A(n8559), .Y(n8330) );
  INVXL U12399 ( .A(n8590), .Y(n8328) );
  AOI2BB2XL U12400 ( .B0(n8434), .B1(n8452), .A0N(n3087), .A1N(n8453), .Y(
        n8602) );
  OAI22XL U12401 ( .A0(n19536), .A1(n3036), .B0(n19542), .B1(n19535), .Y(
        n19806) );
  INVXL U12402 ( .A(n19373), .Y(n19821) );
  INVXL U12403 ( .A(n19392), .Y(n19795) );
  AOI2BB2XL U12404 ( .B0(n3036), .B1(n19543), .A0N(n3036), .A1N(n19535), .Y(
        n19591) );
  INVXL U12405 ( .A(n19389), .Y(n19788) );
  INVXL U12406 ( .A(n19437), .Y(n19902) );
  NOR2XL U12407 ( .A(n23204), .B(n23203), .Y(n19343) );
  AOI2BB2XL U12408 ( .B0(n3041), .B1(n19557), .A0N(n3041), .A1N(n19599), .Y(
        n19661) );
  AOI2BB2XL U12409 ( .B0(n3041), .B1(n19555), .A0N(n3041), .A1N(n19584), .Y(
        n19665) );
  INVXL U12410 ( .A(n19617), .Y(n19666) );
  NAND2XL U12411 ( .A(n3041), .B(n19371), .Y(n19372) );
  NAND2XL U12412 ( .A(n3041), .B(n19445), .Y(n19446) );
  AOI2BB2XL U12413 ( .B0(n3041), .B1(n19426), .A0N(n3041), .A1N(n19928), .Y(
        n19623) );
  AOI2BB2XL U12414 ( .B0(n3041), .B1(n19485), .A0N(n3041), .A1N(n19509), .Y(
        n19617) );
  INVXL U12415 ( .A(n15001), .Y(n15407) );
  NOR2XL U12416 ( .A(n23162), .B(n23161), .Y(n14958) );
  AOI22XL U12417 ( .A0(n3095), .A1(n21662), .B0(n21661), .B1(n21580), .Y(
        n21764) );
  OAI21XL U12418 ( .A0(n14967), .A1(n15221), .B0(n15220), .Y(n15380) );
  NAND2XL U12419 ( .A(n15219), .B(n15256), .Y(n15221) );
  AOI22XL U12420 ( .A0(n15218), .A1(n15355), .B0(n15217), .B1(n15340), .Y(
        n15219) );
  OAI22XL U12421 ( .A0(n15223), .A1(n3101), .B0(n15008), .B1(n15222), .Y(
        n15379) );
  OR2XL U12422 ( .A(n15203), .B(n15359), .Y(n15205) );
  OAI22XL U12423 ( .A0(n15192), .A1(n3101), .B0(n15008), .B1(n15191), .Y(
        n15373) );
  AOI22XL U12424 ( .A0(n3167), .A1(n15246), .B0(n15194), .B1(n15055), .Y(
        n15354) );
  INVXL U12425 ( .A(n23157), .Y(n15038) );
  INVXL U12426 ( .A(n15424), .Y(n15425) );
  OAI22XL U12427 ( .A0(n15153), .A1(n3156), .B0(n3016), .B1(n15152), .Y(n15427) );
  AOI22XL U12428 ( .A0(n15263), .A1(n3034), .B0(n3090), .B1(n15262), .Y(n15432) );
  AOI2BB2XL U12429 ( .B0(n6194), .B1(n15199), .A0N(n6194), .A1N(n15200), .Y(
        n15349) );
  OAI21XL U12430 ( .A0(n21854), .A1(n21789), .B0(n21788), .Y(n21814) );
  AOI22XL U12431 ( .A0(n21785), .A1(n21784), .B0(n21979), .B1(n21803), .Y(
        n21786) );
  OAI21XL U12432 ( .A0(n21854), .A1(n21808), .B0(n21807), .Y(n21818) );
  AOI21XL U12433 ( .A0(n21808), .A1(n3222), .B0(n21849), .Y(n21807) );
  NAND2XL U12434 ( .A(n21806), .B(n21805), .Y(n21808) );
  AOI2BB2XL U12435 ( .B0(n21781), .B1(n3096), .A0N(n3096), .A1N(n21780), .Y(
        n21847) );
  INVXL U12436 ( .A(n21864), .Y(n21865) );
  OAI21XL U12437 ( .A0(n21854), .A1(n21529), .B0(n21528), .Y(n21832) );
  AOI21XL U12438 ( .A0(n21529), .A1(n3222), .B0(n21849), .Y(n21528) );
  OAI211XL U12439 ( .A0(n3171), .A1(n21633), .B0(n21506), .C0(n21526), .Y(
        n21529) );
  NAND2XL U12440 ( .A(n21618), .B(n3171), .Y(n21526) );
  NAND4XL U12441 ( .A(n7894), .B(n7893), .C(n7892), .D(n7891), .Y(n8425) );
  NAND2XL U12442 ( .A(n19346), .B(w2[3]), .Y(n7893) );
  NAND4XL U12443 ( .A(n7899), .B(n7898), .C(n7897), .D(n7896), .Y(n8423) );
  NAND2XL U12444 ( .A(n19346), .B(w2[2]), .Y(n7898) );
  NAND4XL U12445 ( .A(n7929), .B(n7928), .C(n7927), .D(n7926), .Y(n8408) );
  NAND2XL U12446 ( .A(n19346), .B(w2[5]), .Y(n7928) );
  NAND4XL U12447 ( .A(n7924), .B(n7923), .C(n7922), .D(n7921), .Y(n8428) );
  NAND2XL U12448 ( .A(n19346), .B(w2[4]), .Y(n7923) );
  NAND2XL U12449 ( .A(n6217), .B(y10[12]), .Y(n7982) );
  AOI21XL U12450 ( .A0(n23001), .A1(n3218), .B0(n22838), .Y(n22839) );
  OAI2BB1XL U12451 ( .A0N(n11071), .A1N(n22969), .B0(n22970), .Y(n22838) );
  OAI22X1 U12452 ( .A0(n17060), .A1(n16938), .B0(n17061), .B1(n16937), .Y(
        n16974) );
  AOI222XL U12453 ( .A0(n23003), .A1(n11071), .B0(n22969), .B1(n3218), .C0(
        n23001), .C1(n9109), .Y(n22747) );
  INVXL U12454 ( .A(n23021), .Y(n22829) );
  XOR2XL U12455 ( .A(n22668), .B(n3119), .Y(M6_mult_x_15_n1041) );
  INVXL U12456 ( .A(n23143), .Y(M6_mult_x_15_n1018) );
  XOR2XL U12457 ( .A(n22825), .B(n3058), .Y(M6_mult_x_15_n1065) );
  AOI222XL U12458 ( .A0(n22988), .A1(n3219), .B0(n22980), .B1(n11073), .C0(
        n22976), .C1(n11063), .Y(n22785) );
  AOI222XL U12459 ( .A0(n23003), .A1(n3218), .B0(n22969), .B1(n23089), .C0(
        n23001), .C1(n11074), .Y(n22685) );
  XOR2XL U12460 ( .A(n22746), .B(n3056), .Y(M6_mult_x_15_n1087) );
  XNOR2XL U12461 ( .A(n25870), .B(n25872), .Y(n7632) );
  XOR2XL U12462 ( .A(n22916), .B(n3056), .Y(M6_mult_x_15_n1104) );
  XOR2XL U12463 ( .A(n22807), .B(n3221), .Y(M6_mult_x_15_n1201) );
  XNOR2XL U12464 ( .A(n22767), .B(n22766), .Y(n23145) );
  NAND2XL U12465 ( .A(n22765), .B(n22764), .Y(n22766) );
  INVXL U12466 ( .A(n22763), .Y(n22765) );
  XOR2XL U12467 ( .A(n22632), .B(n22631), .Y(n23111) );
  NAND2XL U12468 ( .A(n22630), .B(n22629), .Y(n22631) );
  XNOR2XL U12469 ( .A(n22596), .B(n22595), .Y(n23107) );
  NAND2XL U12470 ( .A(n22594), .B(n22593), .Y(n22595) );
  AOI21XL U12471 ( .A0(n22632), .A1(n22630), .B0(n22591), .Y(n22596) );
  INVXL U12472 ( .A(n22592), .Y(n22594) );
  XOR2XL U12473 ( .A(n22775), .B(n22576), .Y(n23026) );
  NAND2XL U12474 ( .A(n22774), .B(n22772), .Y(n22576) );
  AOI222XL U12475 ( .A0(n22928), .A1(n26496), .B0(n22700), .B1(n10775), .C0(
        n22927), .C1(n10769), .Y(n21076) );
  AOI222XL U12476 ( .A0(n22892), .A1(n23002), .B0(n22708), .B1(n10749), .C0(
        n22891), .C1(n3116), .Y(n22893) );
  AOI222XL U12477 ( .A0(n22988), .A1(n23151), .B0(n22980), .B1(n10789), .C0(
        n22976), .C1(n3220), .Y(n22736) );
  NAND2XL U12478 ( .A(w2[81]), .B(valid[0]), .Y(n11177) );
  NAND2XL U12479 ( .A(w2[49]), .B(n23973), .Y(n11178) );
  XNOR2XL U12480 ( .A(n10751), .B(n10771), .Y(n22978) );
  NAND2XL U12481 ( .A(n10748), .B(n10772), .Y(n10751) );
  INVXL U12482 ( .A(M0_U3_U1_enc_tree_2__2__24_), .Y(M0_U3_U1_or2_inv_2__24_)
         );
  NOR2XL U12483 ( .A(n25870), .B(M0_a_18_), .Y(M0_U3_U1_enc_tree_1__1__12_) );
  INVXL U12484 ( .A(M0_U4_U1_enc_tree_2__2__24_), .Y(M0_U4_U1_or2_inv_2__24_)
         );
  INVXL U12485 ( .A(M0_U4_U1_or2_tree_1__2__24_), .Y(M0_U4_U1_or2_inv_1__24_)
         );
  INVXL U12486 ( .A(M0_U3_U1_or2_tree_1__2__24_), .Y(M0_U3_U1_or2_inv_1__24_)
         );
  OAI22X1 U12487 ( .A0(n6991), .A1(n6286), .B0(n6990), .B1(n6341), .Y(n6343)
         );
  XNOR2XL U12488 ( .A(n4806), .B(n25870), .Y(n6788) );
  XNOR2XL U12489 ( .A(M0_b_1_), .B(n23219), .Y(n6791) );
  XOR2XL U12490 ( .A(n3196), .B(n5718), .Y(n5053) );
  AOI22X1 U12491 ( .A0(n6733), .A1(target_temp[0]), .B0(n4579), .B1(w1[0]), 
        .Y(n6241) );
  AOI22X1 U12492 ( .A0(n6733), .A1(target_temp[4]), .B0(n4579), .B1(w1[4]), 
        .Y(n6269) );
  AOI22X1 U12493 ( .A0(n7389), .A1(target_temp[14]), .B0(n3123), .B1(w1[14]), 
        .Y(n6262) );
  AOI22X1 U12494 ( .A0(n7389), .A1(target_temp[12]), .B0(in_valid_d), .B1(
        w1[12]), .Y(n6249) );
  BUFX3 U12495 ( .A(n6830), .Y(n25876) );
  AOI21X1 U12496 ( .A0(n7389), .A1(y10[12]), .B0(n25150), .Y(n5565) );
  XOR2X1 U12497 ( .A(M3_mult_x_15_b_1_), .B(M3_mult_x_15_b_3_), .Y(n6125) );
  XNOR2XL U12498 ( .A(n18453), .B(M3_mult_x_15_b_13_), .Y(n17551) );
  XOR2X1 U12499 ( .A(n3211), .B(n5957), .Y(n5692) );
  XNOR2XL U12500 ( .A(M3_mult_x_15_b_20_), .B(n17073), .Y(n5067) );
  XNOR2XL U12501 ( .A(n11220), .B(n11219), .Y(n10785) );
  AOI222XL U12502 ( .A0(n22928), .A1(n11059), .B0(n22700), .B1(n11058), .C0(
        n22927), .C1(n23151), .Y(n22791) );
  AOI222XL U12503 ( .A0(n22988), .A1(n11062), .B0(n22980), .B1(n3217), .C0(
        n22976), .C1(n26493), .Y(n22861) );
  AOI222XL U12504 ( .A0(n23003), .A1(n11073), .B0(n22969), .B1(n11063), .C0(
        n23001), .C1(n23109), .Y(n22802) );
  XOR3X2 U12505 ( .A(n16735), .B(n16734), .C(n16733), .Y(n16755) );
  NAND2BXL U12506 ( .AN(n3110), .B(n3022), .Y(n16013) );
  XNOR2X1 U12507 ( .A(M5_mult_x_15_n1), .B(M3_mult_x_15_b_21_), .Y(n16012) );
  XOR2XL U12508 ( .A(n3022), .B(n3208), .Y(n15972) );
  XNOR2X1 U12509 ( .A(M5_mult_x_15_n1), .B(n3202), .Y(n15971) );
  OAI21X2 U12510 ( .A0(n25813), .A1(n26251), .B0(n5019), .Y(n5374) );
  AOI22X1 U12511 ( .A0(n5480), .A1(sigma11[11]), .B0(in_valid_t), .B1(w2[43]), 
        .Y(n5019) );
  INVXL U12512 ( .A(M4_U4_U1_enc_tree_1__1__20_), .Y(M3_U4_U1_or2_inv_1__20_)
         );
  INVXL U12513 ( .A(M3_U4_U1_or2_tree_1__2__24_), .Y(M3_U4_U1_or2_inv_1__24_)
         );
  INVXL U12514 ( .A(M4_U4_U1_enc_tree_1__1__28_), .Y(M3_U4_U1_or2_inv_1__28_)
         );
  INVXL U12515 ( .A(M4_U4_U1_enc_tree_1__1__12_), .Y(M4_U4_U1_or2_inv_1__12_)
         );
  INVXL U12516 ( .A(M4_U4_U1_enc_tree_2__2__24_), .Y(M3_U4_U1_or2_inv_2__24_)
         );
  NOR2XL U12517 ( .A(n25883), .B(M4_a_20_), .Y(M4_U3_U1_enc_tree_1__1__10_) );
  INVXL U12518 ( .A(n22892), .Y(n22709) );
  INVXL U12519 ( .A(n22497), .Y(n22498) );
  INVXL U12520 ( .A(n22496), .Y(n22499) );
  OAI22X1 U12521 ( .A0(n11057), .A1(n26216), .B0(n9107), .B1(n25952), .Y(
        n11160) );
  AOI21XL U12522 ( .A0(n11053), .A1(n11052), .B0(n11051), .Y(n11054) );
  NAND2XL U12523 ( .A(n11048), .B(n11053), .Y(n11055) );
  NAND2XL U12524 ( .A(n11050), .B(n11049), .Y(n11051) );
  NAND2XL U12525 ( .A(n11061), .B(n22601), .Y(n22582) );
  NOR2XL U12526 ( .A(n22575), .B(n22776), .Y(n22586) );
  NOR2XL U12527 ( .A(n22590), .B(n22592), .Y(n11065) );
  AOI21XL U12528 ( .A0(n11065), .A1(n22585), .B0(n11064), .Y(n11066) );
  NAND2XL U12529 ( .A(n22593), .B(n22629), .Y(n11064) );
  AOI21XL U12530 ( .A0(n11061), .A1(n22602), .B0(n11060), .Y(n22584) );
  NAND2XL U12531 ( .A(n22764), .B(n22759), .Y(n11060) );
  OAI22XL U12532 ( .A0(n23193), .A1(n26229), .B0(n9107), .B1(n25940), .Y(
        n11143) );
  AOI21XL U12533 ( .A0(n11076), .A1(n22497), .B0(n11075), .Y(n22504) );
  NAND2XL U12534 ( .A(n22531), .B(n22526), .Y(n11075) );
  NAND2XL U12535 ( .A(n11070), .B(n11072), .Y(n11079) );
  OAI22X1 U12536 ( .A0(n16701), .A1(n16125), .B0(n16699), .B1(n16614), .Y(
        n16162) );
  OAI22XL U12537 ( .A0(n16962), .A1(n16124), .B0(n16960), .B1(n16183), .Y(
        n16163) );
  INVX1 U12538 ( .A(M3_mult_x_15_b_6_), .Y(n16283) );
  OAI22X1 U12539 ( .A0(n16867), .A1(n16312), .B0(n16939), .B1(n16940), .Y(
        n16972) );
  OAI21XL U12540 ( .A0(n19237), .A1(n25941), .B0(n19199), .Y(n19438) );
  NOR2XL U12541 ( .A(n23183), .B(n23182), .Y(n8211) );
  INVXL U12542 ( .A(n8356), .Y(n8402) );
  INVXL U12543 ( .A(n8525), .Y(n8562) );
  NAND2XL U12544 ( .A(n3040), .B(n8480), .Y(n8481) );
  ADDFX2 U12545 ( .A(n6840), .B(n6839), .CI(n6838), .CO(n6914), .S(n6878) );
  OAI22XL U12546 ( .A0(n7633), .A1(n6823), .B0(n6841), .B1(n7634), .Y(n6839)
         );
  OR2X2 U12547 ( .A(n6953), .B(n6952), .Y(n5136) );
  NOR2X1 U12548 ( .A(n19782), .B(n19807), .Y(n19914) );
  OAI22XL U12549 ( .A0(n10541), .A1(n9462), .B0(n10329), .B1(n9506), .Y(n9512)
         );
  OAI21X1 U12550 ( .A0(n9522), .A1(n9523), .B0(n9521), .Y(n5520) );
  XNOR2XL U12551 ( .A(n10494), .B(M2_mult_x_15_n1668), .Y(n10495) );
  INVX1 U12552 ( .A(n10329), .Y(n5758) );
  OAI22XL U12553 ( .A0(n10660), .A1(n10539), .B0(n3178), .B1(n10538), .Y(
        n10513) );
  OAI21XL U12554 ( .A0(n9716), .A1(n9717), .B0(n9715), .Y(n5141) );
  XOR3X2 U12555 ( .A(n9650), .B(n9649), .C(n9648), .Y(n9685) );
  NOR2XL U12556 ( .A(n25885), .B(n5255), .Y(M2_U3_U1_enc_tree_1__1__10_) );
  INVXL U12557 ( .A(M2_U3_U1_enc_tree_0__2__12_), .Y(
        M2_U3_U1_enc_tree_0__3__8_) );
  OAI22XL U12558 ( .A0(n4570), .A1(n9297), .B0(n10403), .B1(n9230), .Y(n9260)
         );
  CMPR32X1 U12559 ( .A(n11726), .B(n11725), .C(n11724), .CO(n11736), .S(n11803) );
  OAI22XL U12560 ( .A0(n12598), .A1(n11673), .B0(n12342), .B1(n11644), .Y(
        n11726) );
  XNOR2XL U12561 ( .A(n12732), .B(n11499), .Y(n11744) );
  XNOR2X1 U12562 ( .A(n12758), .B(n12279), .Y(n11662) );
  OAI22XL U12563 ( .A0(n12717), .A1(n11829), .B0(n12718), .B1(n11745), .Y(
        n11834) );
  XNOR2XL U12564 ( .A(M3_mult_x_15_a_17_), .B(n11499), .Y(n11843) );
  XNOR2XL U12565 ( .A(n12233), .B(n3198), .Y(n11830) );
  XNOR2XL U12566 ( .A(n12271), .B(n12732), .Y(n6115) );
  XNOR2XL U12567 ( .A(n25884), .B(n3197), .Y(n11816) );
  XOR2X1 U12568 ( .A(n25884), .B(n5957), .Y(n5956) );
  XNOR2XL U12569 ( .A(n18638), .B(n3198), .Y(n18544) );
  XOR2X1 U12570 ( .A(n18638), .B(n3208), .Y(n17681) );
  OAI22XL U12571 ( .A0(n18083), .A1(n17870), .B0(n18429), .B1(n17707), .Y(
        n17928) );
  OAI22XL U12572 ( .A0(n13399), .A1(n13721), .B0(n13390), .B1(n13790), .Y(
        n13398) );
  XNOR2XL U12573 ( .A(n14306), .B(n13693), .Y(n13650) );
  XOR2X1 U12574 ( .A(M1_b_2_), .B(M1_b_3_), .Y(n5167) );
  XNOR2XL U12575 ( .A(n14288), .B(n13693), .Y(n13556) );
  OR2XL U12576 ( .A(M1_U4_U1_or2_tree_0__2__16_), .B(
        M1_U4_U1_or2_tree_0__2__24_), .Y(n26212) );
  INVXL U12577 ( .A(M1_U3_U1_enc_tree_0__2__12_), .Y(
        M1_U3_U1_enc_tree_0__3__8_) );
  XNOR2XL U12578 ( .A(n18500), .B(M3_mult_x_15_b_21_), .Y(n17826) );
  XNOR2X1 U12579 ( .A(n18468), .B(n3198), .Y(n17741) );
  XNOR2XL U12580 ( .A(M4_a_17_), .B(n18611), .Y(n17779) );
  XNOR2XL U12581 ( .A(n18638), .B(n18611), .Y(n18545) );
  XNOR2XL U12582 ( .A(n18638), .B(M3_mult_x_15_b_13_), .Y(n17834) );
  OAI22XL U12583 ( .A0(n13934), .A1(n14044), .B0(n13975), .B1(n13974), .Y(
        n13956) );
  OAI22XL U12584 ( .A0(n13933), .A1(n6191), .B0(n13970), .B1(n14298), .Y(
        n13957) );
  CMPR32X1 U12585 ( .A(n13960), .B(n13961), .C(n13959), .CO(n14021), .S(n13954) );
  OAI22XL U12586 ( .A0(n13916), .A1(n14157), .B0(n13962), .B1(n14120), .Y(
        n13959) );
  OAI22XL U12587 ( .A0(n13915), .A1(n14249), .B0(n13963), .B1(n14250), .Y(
        n13960) );
  OAI22XL U12588 ( .A0(n14023), .A1(n14227), .B0(n13963), .B1(n14249), .Y(
        n14018) );
  OAI22XL U12589 ( .A0(n14014), .A1(n14120), .B0(n13962), .B1(n14121), .Y(
        n14019) );
  CMPR32X1 U12590 ( .A(n14013), .B(n14012), .C(n14011), .CO(n14056), .S(n14034) );
  OAI22XL U12591 ( .A0(n13975), .A1(n14044), .B0(n13974), .B1(n14030), .Y(
        n14013) );
  OAI22XL U12592 ( .A0(n14016), .A1(n14198), .B0(n13976), .B1(n14208), .Y(
        n14012) );
  OAI22XL U12593 ( .A0(n14016), .A1(n14208), .B0(n14046), .B1(n14198), .Y(
        n14051) );
  OAI2BB1XL U12594 ( .A0N(n14129), .A1N(n14128), .B0(n14127), .Y(n14141) );
  NAND2XL U12595 ( .A(n14126), .B(n14125), .Y(n14127) );
  XNOR2XL U12596 ( .A(n14265), .B(n23173), .Y(n14189) );
  OAI22XL U12597 ( .A0(n2993), .A1(n14236), .B0(n14289), .B1(n14235), .Y(
        n14194) );
  XNOR2XL U12598 ( .A(n14357), .B(n25862), .Y(n14148) );
  XNOR2X1 U12599 ( .A(n14307), .B(n14228), .Y(n14159) );
  INVXL U12600 ( .A(n14196), .Y(n14152) );
  OAI22XL U12601 ( .A0(n17148), .A1(n3196), .B0(n17147), .B1(n3048), .Y(n17072) );
  XNOR2XL U12602 ( .A(n12732), .B(n3198), .Y(n12638) );
  XOR2X1 U12603 ( .A(n12561), .B(n12732), .Y(n4908) );
  OAI22XL U12604 ( .A0(n18083), .A1(n18082), .B0(n18429), .B1(n6026), .Y(
        n18244) );
  OAI22X1 U12605 ( .A0(n18721), .A1(n12271), .B0(n17512), .B1(
        M3_mult_x_15_b_3_), .Y(n17523) );
  OAI22XL U12606 ( .A0(n17516), .A1(n18429), .B0(n18083), .B1(n5020), .Y(
        n17522) );
  XNOR2XL U12607 ( .A(n14306), .B(n25863), .Y(n14233) );
  XNOR2XL U12608 ( .A(n14357), .B(n25863), .Y(n14252) );
  CLKINVX3 U12609 ( .A(n13428), .Y(n14251) );
  OAI22XL U12610 ( .A0(n2993), .A1(n25864), .B0(n14289), .B1(n14288), .Y(
        n14264) );
  XNOR2XL U12611 ( .A(n14357), .B(n14228), .Y(n14214) );
  OAI22XL U12612 ( .A0(n2993), .A1(n14266), .B0(n14289), .B1(n14265), .Y(
        n14234) );
  OAI22X1 U12613 ( .A0(n13728), .A1(n14120), .B0(n13698), .B1(n14121), .Y(
        n13725) );
  NAND2XL U12614 ( .A(n6053), .B(n3214), .Y(n6050) );
  INVXL U12615 ( .A(n6053), .Y(n6052) );
  INVXL U12616 ( .A(n25864), .Y(n14278) );
  OAI22XL U12617 ( .A0(n14282), .A1(n25863), .B0(n14268), .B1(n14267), .Y(
        n14276) );
  OAI22XL U12618 ( .A0(n2993), .A1(n14288), .B0(n14289), .B1(n14307), .Y(
        n14277) );
  INVXL U12619 ( .A(n23173), .Y(n14290) );
  NAND2X1 U12620 ( .A(in_valid_d), .B(w1[148]), .Y(n11544) );
  OAI22XL U12621 ( .A0(n2993), .A1(n14307), .B0(n14289), .B1(n14306), .Y(
        n14287) );
  NOR2XL U12622 ( .A(n3094), .B(n19665), .Y(n19692) );
  NAND2XL U12623 ( .A(n19415), .B(n19409), .Y(n19417) );
  INVXL U12624 ( .A(n23203), .Y(n19416) );
  NAND2XL U12625 ( .A(n19410), .B(n19415), .Y(n19412) );
  OAI21XL U12626 ( .A0(n3160), .A1(n8348), .B0(n8347), .Y(n8649) );
  AOI21XL U12627 ( .A0(n8348), .A1(n8823), .B0(n3155), .Y(n8347) );
  NAND2XL U12628 ( .A(n8295), .B(n8346), .Y(n8348) );
  AOI21XL U12629 ( .A0(n8711), .A1(n8823), .B0(n3155), .Y(n8710) );
  NAND2XL U12630 ( .A(n8295), .B(n8709), .Y(n8711) );
  NOR2X1 U12631 ( .A(n8654), .B(n3154), .Y(n8785) );
  NAND2XL U12632 ( .A(n8285), .B(n8279), .Y(n8288) );
  INVXL U12633 ( .A(n23178), .Y(n8287) );
  NOR2X1 U12634 ( .A(n8284), .B(n8283), .Y(n8565) );
  AOI22XL U12635 ( .A0(n8592), .A1(n8579), .B0(n3092), .B1(n8562), .Y(n8607)
         );
  NOR2XL U12636 ( .A(n8592), .B(n8572), .Y(n8604) );
  AOI21XL U12637 ( .A0(n19819), .A1(n19952), .B0(n3164), .Y(n19818) );
  NAND2XL U12638 ( .A(n19424), .B(n19817), .Y(n19819) );
  OAI21XL U12639 ( .A0(n3165), .A1(n19793), .B0(n19792), .Y(n19825) );
  AOI21XL U12640 ( .A0(n19793), .A1(n19952), .B0(n3164), .Y(n19792) );
  NAND2XL U12641 ( .A(n19424), .B(n19791), .Y(n19793) );
  AOI22XL U12642 ( .A0(n19790), .A1(n3159), .B0(n19789), .B1(n19807), .Y(
        n19791) );
  OAI21XL U12643 ( .A0(n3165), .A1(n19786), .B0(n19785), .Y(n19823) );
  AOI21XL U12644 ( .A0(n19786), .A1(n19952), .B0(n3164), .Y(n19785) );
  NAND2XL U12645 ( .A(n19424), .B(n19784), .Y(n19786) );
  AOI22XL U12646 ( .A0(n19783), .A1(n3159), .B0(n19782), .B1(n19807), .Y(
        n19784) );
  AOI21XL U12647 ( .A0(n19814), .A1(n19952), .B0(n3164), .Y(n19813) );
  NAND2XL U12648 ( .A(n19424), .B(n19812), .Y(n19814) );
  AOI21XL U12649 ( .A0(n19900), .A1(n19952), .B0(n3164), .Y(n19899) );
  NAND2XL U12650 ( .A(n19424), .B(n19898), .Y(n19900) );
  INVXL U12651 ( .A(n19903), .Y(n19982) );
  NOR2XL U12652 ( .A(n23163), .B(n23164), .Y(n14959) );
  NOR2XL U12653 ( .A(n23160), .B(n23159), .Y(n14961) );
  AOI22XL U12654 ( .A0(n15333), .A1(n15324), .B0(n15337), .B1(n15323), .Y(
        n15331) );
  NOR4BXL U12655 ( .AN(n15311), .B(n15310), .C(n15309), .D(n15308), .Y(n15344)
         );
  NAND2XL U12656 ( .A(n3016), .B(n15055), .Y(n15295) );
  OAI21XL U12657 ( .A0(n21854), .A1(n21655), .B0(n21654), .Y(n21759) );
  NAND2XL U12658 ( .A(n21805), .B(n21653), .Y(n21655) );
  OAI21XL U12659 ( .A0(n21854), .A1(n21638), .B0(n21637), .Y(n21757) );
  NAND2XL U12660 ( .A(n21805), .B(n21636), .Y(n21638) );
  INVXL U12661 ( .A(n21620), .Y(n21657) );
  INVXL U12662 ( .A(n23119), .Y(n21493) );
  NAND2XL U12663 ( .A(n21256), .B(w1[22]), .Y(n21310) );
  NAND2XL U12664 ( .A(n21256), .B(w1[18]), .Y(n21299) );
  INVXL U12665 ( .A(n21775), .Y(n21195) );
  NOR2XL U12666 ( .A(n15380), .B(n15379), .Y(n15643) );
  NAND2XL U12667 ( .A(n15380), .B(n15379), .Y(n15644) );
  NOR2XL U12668 ( .A(n15602), .B(n15606), .Y(n15609) );
  INVXL U12669 ( .A(n15601), .Y(n15602) );
  AOI21XL U12670 ( .A0(n15682), .A1(n15390), .B0(n15389), .Y(n15391) );
  INVXL U12671 ( .A(n15681), .Y(n15389) );
  INVXL U12672 ( .A(n15675), .Y(n15390) );
  OAI21XL U12673 ( .A0(n21854), .A1(n21577), .B0(n21576), .Y(n21824) );
  AOI21XL U12674 ( .A0(n21577), .A1(n3222), .B0(n21849), .Y(n21576) );
  AOI22XL U12675 ( .A0(n21574), .A1(n21573), .B0(n21803), .B1(n21994), .Y(
        n21575) );
  OAI21XL U12676 ( .A0(n21854), .A1(n21615), .B0(n21614), .Y(n21822) );
  AOI21XL U12677 ( .A0(n21615), .A1(n3222), .B0(n21849), .Y(n21614) );
  NAND2XL U12678 ( .A(n21613), .B(n21805), .Y(n21615) );
  AOI22XL U12679 ( .A0(n21612), .A1(n21803), .B0(n21611), .B1(n21801), .Y(
        n21613) );
  NAND2XL U12680 ( .A(n21814), .B(n21813), .Y(n22086) );
  NOR2XL U12681 ( .A(n21818), .B(n21817), .Y(n22080) );
  AOI21XL U12682 ( .A0(n21792), .A1(n21816), .B0(n21815), .Y(n22078) );
  INVXL U12683 ( .A(n22086), .Y(n21815) );
  INVXL U12684 ( .A(n22089), .Y(n21816) );
  NAND2XL U12685 ( .A(n22090), .B(n21792), .Y(n22079) );
  NAND2XL U12686 ( .A(n21818), .B(n21817), .Y(n22081) );
  INVXL U12687 ( .A(n21509), .Y(n21993) );
  INVXL U12688 ( .A(n21511), .Y(n21998) );
  NOR2XL U12689 ( .A(n22079), .B(n22080), .Y(n21820) );
  OAI21XL U12690 ( .A0(n22078), .A1(n22080), .B0(n22081), .Y(n21819) );
  NAND2XL U12691 ( .A(n21832), .B(n21831), .Y(n22107) );
  OAI21XL U12692 ( .A0(n21830), .A1(n22113), .B0(n21829), .Y(n22104) );
  INVXL U12693 ( .A(n22112), .Y(n21828) );
  INVXL U12694 ( .A(n22118), .Y(n21827) );
  OAI21XL U12695 ( .A0(n21854), .A1(n21861), .B0(n21860), .Y(n21887) );
  AOI21XL U12696 ( .A0(n21861), .A1(n3222), .B0(n21849), .Y(n21860) );
  OAI211XL U12697 ( .A0(n3171), .A1(n21858), .B0(n21506), .C0(n21857), .Y(
        n21861) );
  OAI22XL U12698 ( .A0(n17074), .A1(n17073), .B0(n16319), .B1(n3212), .Y(
        n17081) );
  OAI22XL U12699 ( .A0(n17148), .A1(n3048), .B0(n17147), .B1(
        M3_mult_x_15_b_20_), .Y(n17082) );
  OAI22X1 U12700 ( .A0(n12715), .A1(n11663), .B0(n12525), .B1(n11629), .Y(
        n11666) );
  OAI22X1 U12701 ( .A0(n12618), .A1(n11651), .B0(n12119), .B1(n11641), .Y(
        n11669) );
  XNOR2X1 U12702 ( .A(n3211), .B(n3048), .Y(n16959) );
  CMPR32X1 U12703 ( .A(n16958), .B(n16957), .C(n16956), .CO(n16999), .S(n17019) );
  OAI22XL U12704 ( .A0(n17074), .A1(n16320), .B0(n16319), .B1(n16981), .Y(
        n16956) );
  OAI22XL U12705 ( .A0(n12598), .A1(n11644), .B0(n12342), .B1(n11655), .Y(
        n11661) );
  NAND2X1 U12706 ( .A(n5594), .B(n5593), .Y(n7666) );
  OAI21XL U12707 ( .A0(n7576), .A1(n7577), .B0(n7575), .Y(n5594) );
  NAND2XL U12708 ( .A(n9105), .B(n9104), .Y(n11209) );
  NAND2XL U12709 ( .A(w2[72]), .B(valid[0]), .Y(n9104) );
  NAND2XL U12710 ( .A(w2[40]), .B(n23973), .Y(n9105) );
  INVXL U12711 ( .A(n23149), .Y(M6_mult_x_15_n1020) );
  XOR2XL U12712 ( .A(n22885), .B(n3119), .Y(M6_mult_x_15_n1043) );
  XOR2XL U12713 ( .A(n22890), .B(n3054), .Y(M6_mult_x_15_n1139) );
  XOR2XL U12714 ( .A(n22854), .B(n3058), .Y(M6_mult_x_15_n1067) );
  XOR2XL U12715 ( .A(n22574), .B(n3056), .Y(M6_mult_x_15_n1086) );
  XOR2XL U12716 ( .A(n22600), .B(n3055), .Y(M6_mult_x_15_n1110) );
  XOR2XL U12717 ( .A(n21066), .B(n3056), .Y(M6_mult_x_15_n1084) );
  XOR2XL U12718 ( .A(n22561), .B(n3119), .Y(M6_mult_x_15_n1036) );
  INVXL U12719 ( .A(n23112), .Y(M6_mult_x_15_n1013) );
  XOR2XL U12720 ( .A(n22566), .B(n3056), .Y(M6_mult_x_15_n1085) );
  INVXL U12721 ( .A(n23136), .Y(M6_mult_x_15_n1014) );
  XOR2XL U12722 ( .A(n22666), .B(n3221), .Y(M6_mult_x_15_n1198) );
  XOR2XL U12723 ( .A(n22688), .B(n3221), .Y(M6_mult_x_15_n1196) );
  XOR2XL U12724 ( .A(n22809), .B(n3056), .Y(M6_mult_x_15_n1100) );
  XOR2XL U12725 ( .A(n22873), .B(n3053), .Y(M6_mult_x_15_n1172) );
  XOR2XL U12726 ( .A(n22516), .B(n22508), .Y(n23091) );
  NAND2XL U12727 ( .A(n11070), .B(n22507), .Y(n22508) );
  INVXL U12728 ( .A(n22507), .Y(n22515) );
  NAND2XL U12729 ( .A(n11071), .B(n3218), .Y(n22517) );
  INVXL U12730 ( .A(n22943), .Y(n22960) );
  INVXL U12731 ( .A(M6_mult_x_15_n634), .Y(n22961) );
  AOI222XL U12732 ( .A0(n22892), .A1(n10769), .B0(n22708), .B1(n23002), .C0(
        n22891), .C1(n10749), .Y(n22857) );
  AOI222XL U12733 ( .A0(n22988), .A1(n11058), .B0(n22980), .B1(n23151), .C0(
        n22976), .C1(n10789), .Y(n22677) );
  AOI222XL U12734 ( .A0(n22928), .A1(n10789), .B0(n22700), .B1(n3220), .C0(
        n22927), .C1(n26496), .Y(n22816) );
  AOI21XL U12735 ( .A0(n22952), .A1(n3218), .B0(n22898), .Y(n22899) );
  OAI2BB1XL U12736 ( .A0N(n11071), .A1N(n22897), .B0(n22896), .Y(n22898) );
  AOI222XL U12737 ( .A0(n23023), .A1(n11073), .B0(n22887), .B1(n11063), .C0(
        n23021), .C1(n23109), .Y(n22818) );
  XOR2XL U12738 ( .A(n22866), .B(n21089), .Y(M6_mult_x_15_n1121) );
  NAND3XL U12739 ( .A(n26195), .B(y11[0]), .C(n23973), .Y(n10750) );
  NAND3XL U12740 ( .A(n26195), .B(y11[1]), .C(n23973), .Y(n10746) );
  BUFX3 U12741 ( .A(M0_b_21_), .Y(n7800) );
  BUFX3 U12742 ( .A(M0_b_20_), .Y(n25873) );
  NAND2X1 U12743 ( .A(n5604), .B(w2[22]), .Y(n5607) );
  OAI21XL U12744 ( .A0(n6274), .A1(n26231), .B0(n6273), .Y(n6828) );
  OAI21X1 U12745 ( .A0(n5626), .A1(n5625), .B0(n5624), .Y(n6710) );
  AOI21X1 U12746 ( .A0(n6671), .A1(n5553), .B0(n6670), .Y(n5550) );
  XOR3X2 U12747 ( .A(n6698), .B(n6697), .C(n6699), .Y(n6703) );
  NAND2X1 U12748 ( .A(n5618), .B(n5617), .Y(n6692) );
  NAND2XL U12749 ( .A(n6533), .B(n6532), .Y(n5617) );
  OAI22XL U12750 ( .A0(n6283), .A1(n7512), .B0(n7511), .B1(n6287), .Y(n6358)
         );
  OAI21XL U12751 ( .A0(n7094), .A1(n5131), .B0(n5130), .Y(n6818) );
  ADDFX2 U12752 ( .A(n6773), .B(n6772), .CI(n6771), .CO(n6877), .S(n6766) );
  OAI22XL U12753 ( .A0(n17148), .A1(M3_mult_x_15_b_20_), .B0(n17147), .B1(
        M3_mult_x_15_b_21_), .Y(n17091) );
  OAI22XL U12754 ( .A0(n17060), .A1(n16876), .B0(n17061), .B1(n16870), .Y(
        n16882) );
  OAI21XL U12755 ( .A0(n16962), .A1(n5947), .B0(n5944), .Y(n16879) );
  INVXL U12756 ( .A(M3_U3_U1_or2_tree_0__2__24_), .Y(M3_U3_U1_or2_inv_0__24_)
         );
  XOR2XL U12757 ( .A(n22875), .B(n3119), .Y(M6_mult_x_15_n1045) );
  XOR2XL U12758 ( .A(n22784), .B(n3053), .Y(M6_mult_x_15_n1165) );
  XOR2XL U12759 ( .A(n22920), .B(n3055), .Y(M6_mult_x_15_n1117) );
  XOR2XL U12760 ( .A(n22788), .B(n3058), .Y(M6_mult_x_15_n1071) );
  XOR2XL U12761 ( .A(n22758), .B(n3119), .Y(M6_mult_x_15_n1047) );
  XOR2XL U12762 ( .A(n22835), .B(n11220), .Y(M6_mult_x_15_n1191) );
  XOR2XL U12763 ( .A(n22842), .B(n3056), .Y(M6_mult_x_15_n1095) );
  XNOR2XL U12764 ( .A(n25883), .B(M3_mult_x_15_b_21_), .Y(n18635) );
  XNOR2XL U12765 ( .A(n25883), .B(n3202), .Y(n18651) );
  NOR2X1 U12766 ( .A(n16755), .B(n16754), .Y(n16758) );
  INVX1 U12767 ( .A(n16416), .Y(n5855) );
  OAI22XL U12768 ( .A0(n17288), .A1(n17266), .B0(M3_U4_U1_enc_tree_1__4__16_), 
        .B1(M5_U3_U1_enc_tree_1__4__16_), .Y(n17286) );
  NOR2XL U12769 ( .A(n18822), .B(n17287), .Y(n17266) );
  AOI22X1 U12770 ( .A0(n5480), .A1(sigma11[3]), .B0(in_valid_t), .B1(w2[35]), 
        .Y(n5882) );
  NAND2X1 U12771 ( .A(n5480), .B(sigma11[7]), .Y(n6090) );
  AOI22X1 U12772 ( .A0(n5480), .A1(target_temp[13]), .B0(in_valid_t), .B1(
        learning_rate[13]), .Y(n11490) );
  NAND2X1 U12773 ( .A(n5480), .B(target_temp[9]), .Y(n6163) );
  INVXL U12774 ( .A(n18818), .Y(n18797) );
  NAND2XL U12775 ( .A(n12944), .B(M4_U4_U1_enc_tree_3__3__24_), .Y(n18800) );
  INVXL U12776 ( .A(M4_U4_U1_enc_tree_3__3__16_), .Y(n12944) );
  AND2XL U12777 ( .A(M4_U3_U1_enc_tree_1__1__12_), .B(
        M4_U3_U1_enc_tree_1__1__14_), .Y(n25985) );
  OR2XL U12778 ( .A(M4_U3_U1_enc_tree_2__2__16_), .B(
        M4_U3_U1_enc_tree_2__2__24_), .Y(n26200) );
  XNOR2XL U12779 ( .A(n22534), .B(n22533), .Y(n23098) );
  NAND2XL U12780 ( .A(n22532), .B(n22531), .Y(n22533) );
  AOI21XL U12781 ( .A0(n22529), .A1(n22528), .B0(n22527), .Y(n22534) );
  INVXL U12782 ( .A(n22530), .Y(n22532) );
  NOR2XL U12783 ( .A(n11340), .B(n11042), .Y(n10942) );
  OAI2BB1XL U12784 ( .A0N(n5835), .A1N(n16704), .B0(n3047), .Y(n16180) );
  OAI22XL U12785 ( .A0(n16167), .A1(n3105), .B0(n16977), .B1(n5037), .Y(n16182) );
  XOR2XL U12786 ( .A(n3199), .B(n5718), .Y(n16313) );
  INVXL U12787 ( .A(n9015), .Y(n20445) );
  OAI22XL U12788 ( .A0(n4642), .A1(n7696), .B0(n7712), .B1(n23219), .Y(n7710)
         );
  INVX1 U12789 ( .A(n10316), .Y(n5222) );
  NOR2X1 U12790 ( .A(n10317), .B(n10318), .Y(n5223) );
  NAND2XL U12791 ( .A(n9569), .B(n9568), .Y(n5224) );
  OAI22XL U12792 ( .A0(n10660), .A1(n10515), .B0(n10659), .B1(
        M2_mult_x_15_n1669), .Y(n10537) );
  INVXL U12793 ( .A(n10539), .Y(n10527) );
  OAI22XL U12794 ( .A0(n10517), .A1(n10494), .B0(n10533), .B1(n5079), .Y(
        n10525) );
  OAI22XL U12795 ( .A0(n10660), .A1(n10538), .B0(n10659), .B1(n10515), .Y(
        n10526) );
  INVXL U12796 ( .A(n10585), .Y(n10588) );
  AND2XL U12797 ( .A(n10005), .B(n10004), .Y(n10009) );
  NAND2X1 U12798 ( .A(n5744), .B(n5743), .Y(n10047) );
  OAI21XL U12799 ( .A0(n9830), .A1(n9831), .B0(n5745), .Y(n5744) );
  OAI2BB1X1 U12800 ( .A0N(n9789), .A1N(n9788), .B0(n5765), .Y(n9828) );
  OAI21XL U12801 ( .A0(n9788), .A1(n9789), .B0(n9787), .Y(n5765) );
  XOR2X1 U12802 ( .A(n9823), .B(n5285), .Y(n10014) );
  NOR2X1 U12803 ( .A(n5176), .B(n10044), .Y(n10046) );
  OAI2BB1XL U12804 ( .A0N(n11887), .A1N(n11886), .B0(n11885), .Y(n11905) );
  NAND2XL U12805 ( .A(n11884), .B(n11883), .Y(n11885) );
  OAI22XL U12806 ( .A0(n12715), .A1(n12524), .B0(n12746), .B1(n12514), .Y(
        n12528) );
  OAI22X1 U12807 ( .A0(n12635), .A1(n4890), .B0(n12519), .B1(n12513), .Y(
        n12532) );
  OAI22XL U12808 ( .A0(n12535), .A1(n12701), .B0(n12995), .B1(n3198), .Y(
        n12559) );
  OAI22XL U12809 ( .A0(n12535), .A1(n18673), .B0(n12995), .B1(
        M3_mult_x_15_b_21_), .Y(n12750) );
  XNOR2XL U12810 ( .A(n12751), .B(n5718), .Y(n12700) );
  XNOR2XL U12811 ( .A(n12732), .B(n3202), .Y(n12714) );
  OAI22XL U12812 ( .A0(n12535), .A1(n3196), .B0(n12995), .B1(n3048), .Y(n12730) );
  OAI22X1 U12813 ( .A0(n18433), .A1(n18541), .B0(n5893), .B1(n18453), .Y(
        n18436) );
  OAI22XL U12814 ( .A0(n12715), .A1(n12732), .B0(n12746), .B1(n12731), .Y(
        n12740) );
  OAI22XL U12815 ( .A0(n12535), .A1(n3048), .B0(n12995), .B1(n18673), .Y(
        n12741) );
  NOR2X1 U12816 ( .A(n18520), .B(n18483), .Y(n5445) );
  ADDFX2 U12817 ( .A(n5430), .B(M3_mult_x_15_b_9_), .CI(n18523), .CO(n18549), 
        .S(n18552) );
  OAI21XL U12818 ( .A0(n17952), .A1(n17951), .B0(n17950), .Y(n4834) );
  OAI21X1 U12819 ( .A0(n18624), .A1(n17601), .B0(n5897), .Y(n17660) );
  OAI22XL U12820 ( .A0(n18107), .A1(n17603), .B0(n17902), .B1(n17581), .Y(
        n17661) );
  INVX1 U12821 ( .A(n13347), .Y(n5024) );
  OAI22XL U12822 ( .A0(n13677), .A1(n14298), .B0(n13603), .B1(n6191), .Y(
        n13664) );
  CMPR32X1 U12823 ( .A(n13630), .B(n13629), .C(n13628), .CO(n13710), .S(n13610) );
  OAI22XL U12824 ( .A0(n13568), .A1(n14249), .B0(n13616), .B1(n14250), .Y(
        n13628) );
  OAI22XL U12825 ( .A0(n13567), .A1(n6191), .B0(n13603), .B1(n14298), .Y(
        n13629) );
  OAI22X1 U12826 ( .A0(n18522), .A1(n17741), .B0(n3195), .B1(n17790), .Y(n4885) );
  OAI22XL U12827 ( .A0(n18541), .A1(n17749), .B0(n18539), .B1(n17784), .Y(
        n17775) );
  OAI22XL U12828 ( .A0(n12717), .A1(n11877), .B0(n12718), .B1(n11916), .Y(
        n11924) );
  CMPR32X1 U12829 ( .A(n12614), .B(n12613), .C(n12612), .CO(n12656), .S(n12677) );
  OAI22XL U12830 ( .A0(n12715), .A1(n11985), .B0(n12746), .B1(n12639), .Y(
        n12612) );
  ADDFX2 U12831 ( .A(n12624), .B(n12623), .CI(n12622), .CO(n12654), .S(n12676)
         );
  OAI22X1 U12832 ( .A0(n18659), .A1(n17527), .B0(n17832), .B1(n17554), .Y(
        n17543) );
  OAI22XL U12833 ( .A0(n18541), .A1(n17535), .B0(n5893), .B1(n17552), .Y(
        n17544) );
  AND2X1 U12834 ( .A(n17541), .B(n17540), .Y(n17584) );
  XNOR2XL U12835 ( .A(n18638), .B(n3202), .Y(n18623) );
  XNOR3X2 U12836 ( .A(n5870), .B(n17626), .C(n17625), .Y(n17645) );
  NAND2X1 U12837 ( .A(n17609), .B(n3169), .Y(n5476) );
  INVX1 U12838 ( .A(M3_mult_x_15_b_20_), .Y(n5960) );
  OAI22XL U12839 ( .A0(n18721), .A1(n18673), .B0(n17512), .B1(
        M3_mult_x_15_b_21_), .Y(n18657) );
  NAND3X1 U12840 ( .A(n14663), .B(n23588), .C(n23481), .Y(n14664) );
  NOR2XL U12841 ( .A(n20157), .B(n20175), .Y(n20158) );
  NAND4XL U12842 ( .A(n20177), .B(n20156), .C(n20204), .D(n20203), .Y(n20157)
         );
  NAND2XL U12843 ( .A(n8461), .B(n8898), .Y(n8899) );
  NAND2XL U12844 ( .A(n8894), .B(n8893), .Y(n8895) );
  OAI21XL U12845 ( .A0(n8904), .A1(n8891), .B0(n8890), .Y(n8896) );
  INVXL U12846 ( .A(n8892), .Y(n8894) );
  NAND2XL U12847 ( .A(n8902), .B(n8901), .Y(n8903) );
  INVXL U12848 ( .A(n8732), .Y(n8746) );
  NAND2XL U12849 ( .A(n8706), .B(n8705), .Y(n8724) );
  INVXL U12850 ( .A(n8917), .Y(n8760) );
  NOR2XL U12851 ( .A(n8759), .B(n8919), .Y(n8762) );
  INVXL U12852 ( .A(n8918), .Y(n8759) );
  NAND2XL U12853 ( .A(n8715), .B(n8714), .Y(n8855) );
  AOI21XL U12854 ( .A0(n8797), .A1(n8823), .B0(n3155), .Y(n8796) );
  NAND2XL U12855 ( .A(n8704), .B(n8703), .Y(n8728) );
  NAND2XL U12856 ( .A(n8403), .B(n8931), .Y(n8932) );
  INVXL U12857 ( .A(n19874), .Y(n19862) );
  NAND2XL U12858 ( .A(n19870), .B(n19875), .Y(n19864) );
  AOI21XL U12859 ( .A0(n19989), .A1(n19858), .B0(n19849), .Y(n19850) );
  INVXL U12860 ( .A(n19857), .Y(n19849) );
  NAND2XL U12861 ( .A(n19982), .B(n19858), .Y(n19851) );
  INVXL U12862 ( .A(n19848), .Y(n19858) );
  INVXL U12863 ( .A(n19861), .Y(n19875) );
  INVXL U12864 ( .A(n19871), .Y(n19872) );
  INVXL U12865 ( .A(n20177), .Y(n20201) );
  INVXL U12866 ( .A(n20005), .Y(n20006) );
  NAND2XL U12867 ( .A(n20004), .B(n20007), .Y(n20010) );
  AOI21XL U12868 ( .A0(n19989), .A1(n19988), .B0(n19987), .Y(n19990) );
  INVXL U12869 ( .A(n19983), .Y(n19986) );
  NAND2XL U12870 ( .A(n19982), .B(n19988), .Y(n19991) );
  NAND2XL U12871 ( .A(n19905), .B(n19904), .Y(n19994) );
  NAND2XL U12872 ( .A(n19982), .B(n19980), .Y(n19837) );
  NAND2XL U12873 ( .A(n19844), .B(n19843), .Y(n19984) );
  NAND2XL U12874 ( .A(n19534), .B(n20060), .Y(n20061) );
  NAND2XL U12875 ( .A(n20050), .B(n20049), .Y(n20051) );
  INVXL U12876 ( .A(n20048), .Y(n20050) );
  INVXL U12877 ( .A(n20188), .Y(n20218) );
  INVXL U12878 ( .A(n15823), .Y(n15806) );
  INVXL U12879 ( .A(n15481), .Y(n15495) );
  INVXL U12880 ( .A(n15801), .Y(n15830) );
  INVXL U12881 ( .A(n15809), .Y(n15831) );
  NAND2XL U12882 ( .A(n21759), .B(n21758), .Y(n22095) );
  INVXL U12883 ( .A(n22126), .Y(n22094) );
  OAI21XL U12884 ( .A0(n21854), .A1(n21774), .B0(n21773), .Y(n21812) );
  AOI22XL U12885 ( .A0(n21771), .A1(n21770), .B0(n21974), .B1(n21803), .Y(
        n21772) );
  NOR2XL U12886 ( .A(n21812), .B(n21811), .Y(n22085) );
  OAI21XL U12887 ( .A0(n21762), .A1(n22093), .B0(n21761), .Y(n22077) );
  NAND2XL U12888 ( .A(n22127), .B(n6216), .Y(n21762) );
  AOI21XL U12889 ( .A0(n6216), .A1(n22094), .B0(n21760), .Y(n21761) );
  INVXL U12890 ( .A(n22095), .Y(n21760) );
  NAND2XL U12891 ( .A(n21757), .B(n21756), .Y(n22126) );
  OR2XL U12892 ( .A(n21854), .B(n21668), .Y(n21669) );
  AOI22XL U12893 ( .A0(n21803), .A1(n21872), .B0(n21667), .B1(n21666), .Y(
        n21668) );
  OAI21XL U12894 ( .A0(n21468), .A1(n21478), .B0(n21480), .Y(n21449) );
  INVXL U12895 ( .A(n21481), .Y(n21447) );
  NAND2XL U12896 ( .A(n23394), .B(n21486), .Y(n21487) );
  INVXL U12897 ( .A(n21461), .Y(n21881) );
  INVXL U12898 ( .A(n21520), .Y(n21983) );
  NAND2XL U12899 ( .A(n21311), .B(temp0[18]), .Y(n21300) );
  INVXL U12900 ( .A(n15172), .Y(n15191) );
  INVXL U12901 ( .A(n15226), .Y(n15242) );
  INVXL U12902 ( .A(n15228), .Y(n15259) );
  NAND2XL U12903 ( .A(n15386), .B(n15385), .Y(n15675) );
  INVXL U12904 ( .A(n15674), .Y(n15665) );
  NAND2XL U12905 ( .A(n21824), .B(n21823), .Y(n22112) );
  NAND2XL U12906 ( .A(n21822), .B(n21821), .Y(n22113) );
  INVXL U12907 ( .A(n22111), .Y(n22102) );
  AOI21XL U12908 ( .A0(n21755), .A1(n3222), .B0(n21849), .Y(n21754) );
  NAND2XL U12909 ( .A(n8912), .B(n8925), .Y(n8913) );
  INVXL U12910 ( .A(n8926), .Y(n8911) );
  NAND2XL U12911 ( .A(n8915), .B(n8926), .Y(n8916) );
  AOI21XL U12912 ( .A0(n8131), .A1(n8130), .B0(n8129), .Y(n8132) );
  NAND2X1 U12913 ( .A(n5081), .B(n17132), .Y(n17372) );
  ADDFX2 U12914 ( .A(n17080), .B(n17079), .CI(n17078), .CO(n17135), .S(n17129)
         );
  INVX1 U12915 ( .A(n11755), .Y(n4864) );
  NOR2XL U12916 ( .A(M6_mult_x_15_n528), .B(M6_mult_x_15_n537), .Y(n11028) );
  NAND2XL U12917 ( .A(M6_mult_x_15_n509), .B(M6_mult_x_15_n517), .Y(n11096) );
  XNOR3X2 U12918 ( .A(n7575), .B(n5595), .C(n7576), .Y(n7663) );
  NOR2XL U12919 ( .A(M6_mult_x_15_n491), .B(M6_mult_x_15_n499), .Y(n11036) );
  NAND2XL U12920 ( .A(M6_mult_x_15_n491), .B(M6_mult_x_15_n499), .Y(n11354) );
  NOR2XL U12921 ( .A(n11101), .B(n11114), .Y(n11038) );
  NOR2XL U12922 ( .A(M6_mult_x_15_n549), .B(M6_mult_x_15_n559), .Y(n11042) );
  INVXL U12923 ( .A(n11030), .Y(n11348) );
  XOR2XL U12924 ( .A(n22514), .B(n3119), .Y(M6_mult_x_15_n1035) );
  XOR2XL U12925 ( .A(n22521), .B(n3058), .Y(M6_mult_x_15_n1059) );
  NAND2XL U12926 ( .A(M6_mult_x_15_n626), .B(M6_mult_x_15_n636), .Y(n10931) );
  NAND2XL U12927 ( .A(M6_mult_x_15_n637), .B(M6_mult_x_15_n646), .Y(n10932) );
  NOR2XL U12928 ( .A(M6_mult_x_15_n626), .B(M6_mult_x_15_n636), .Y(n10933) );
  NOR2XL U12929 ( .A(M6_mult_x_15_n637), .B(M6_mult_x_15_n646), .Y(n10744) );
  NAND2XL U12930 ( .A(n10927), .B(n10745), .Y(n10930) );
  OR2XL U12931 ( .A(M6_mult_x_15_n657), .B(M6_mult_x_15_n666), .Y(n10745) );
  AOI21XL U12932 ( .A0(n10927), .A1(n10926), .B0(n10925), .Y(n10928) );
  AND2XL U12933 ( .A(M6_mult_x_15_n647), .B(M6_mult_x_15_n656), .Y(n10925) );
  AOI21XL U12934 ( .A0(n10924), .A1(n10923), .B0(n10922), .Y(n10929) );
  XOR2XL U12935 ( .A(n22902), .B(n3053), .Y(M6_mult_x_15_n1171) );
  XOR2XL U12936 ( .A(n22860), .B(n3054), .Y(M6_mult_x_15_n1147) );
  XNOR2XL U12937 ( .A(n22519), .B(n22518), .Y(n23095) );
  NAND2XL U12938 ( .A(n11072), .B(n22517), .Y(n22518) );
  AOI21XL U12939 ( .A0(n22516), .A1(n11070), .B0(n22515), .Y(n22519) );
  XOR2XL U12940 ( .A(n22771), .B(n3053), .Y(M6_mult_x_15_n1170) );
  XOR2XL U12941 ( .A(n22805), .B(n21089), .Y(M6_mult_x_15_n1122) );
  INVXL U12942 ( .A(n11259), .Y(n11275) );
  INVXL U12943 ( .A(M0_U4_U1_enc_tree_0__4__16_), .Y(n10731) );
  INVXL U12944 ( .A(M0_U4_U1_enc_tree_0__2__12_), .Y(
        M0_U4_U1_enc_tree_0__3__8_) );
  INVXL U12945 ( .A(M0_U3_U1_enc_tree_0__4__16_), .Y(n10730) );
  INVXL U12946 ( .A(M0_U3_U1_enc_tree_0__2__12_), .Y(
        M0_U3_U1_enc_tree_0__3__8_) );
  INVXL U12947 ( .A(n17566), .Y(n5907) );
  OAI22XL U12948 ( .A0(n17060), .A1(n16923), .B0(n17061), .B1(n17039), .Y(
        n17037) );
  NAND2XL U12949 ( .A(M6_mult_x_15_n549), .B(M6_mult_x_15_n559), .Y(n11336) );
  OAI22XL U12950 ( .A0(n18652), .A1(n18638), .B0(n18653), .B1(n18637), .Y(
        n18646) );
  OAI22XL U12951 ( .A0(n18721), .A1(n3048), .B0(n17512), .B1(n18673), .Y(
        n18647) );
  INVXL U12952 ( .A(M5_U3_U1_or2_tree_0__2__24_), .Y(M5_U3_U1_or2_inv_0__24_)
         );
  AOI21XL U12953 ( .A0(n4796), .A1(n5646), .B0(M5_a_12_), .Y(
        M5_U3_U1_enc_tree_0__1__18_) );
  OR2XL U12954 ( .A(M5_U3_U1_or2_tree_0__2__16_), .B(
        M5_U3_U1_or2_tree_0__2__24_), .Y(n26208) );
  NOR2XL U12955 ( .A(n3199), .B(n3211), .Y(M5_U3_U1_or2_tree_0__1__16_) );
  AOI22X1 U12956 ( .A0(n5770), .A1(data[68]), .B0(w2[36]), .B1(in_valid_t), 
        .Y(n5375) );
  INVXL U12957 ( .A(n5470), .Y(n5471) );
  NAND2X1 U12958 ( .A(n5015), .B(data[82]), .Y(n5014) );
  NOR2X2 U12959 ( .A(n4860), .B(n4726), .Y(n5469) );
  AND2X2 U12960 ( .A(in_valid_t), .B(w2[45]), .Y(n4659) );
  NOR2X1 U12961 ( .A(n4860), .B(n26443), .Y(n5468) );
  NOR2BXL U12962 ( .AN(n18428), .B(M4_a_9_), .Y(M4_U3_U1_or2_tree_0__1__20_)
         );
  INVXL U12963 ( .A(M4_U4_U1_or2_tree_0__1__28_), .Y(M3_U4_U1_or2_inv_0__28_)
         );
  INVXL U12964 ( .A(M3_mult_x_15_b_13_), .Y(M3_U4_U1_or2_inv_0__18_) );
  INVXL U12965 ( .A(M4_U3_U1_enc_tree_3__3__16_), .Y(n18798) );
  NOR2XL U12966 ( .A(n21067), .B(n11071), .Y(n11080) );
  INVXL U12967 ( .A(n21068), .Y(n11081) );
  XNOR2XL U12968 ( .A(n21069), .B(n11071), .Y(n23076) );
  AOI21XL U12969 ( .A0(n22570), .A1(n21068), .B0(n21067), .Y(n21069) );
  INVXL U12970 ( .A(n10999), .Y(n10949) );
  INVXL U12971 ( .A(n11350), .Y(n10950) );
  NOR2XL U12972 ( .A(n11006), .B(n11020), .Y(n11024) );
  NOR2XL U12973 ( .A(n11028), .B(n11031), .Y(n10986) );
  NOR2XL U12974 ( .A(n10990), .B(n10992), .Y(n10944) );
  INVXL U12975 ( .A(n20415), .Y(n20463) );
  NOR2XL U12976 ( .A(n3124), .B(n20434), .Y(n20412) );
  INVXL U12977 ( .A(n20461), .Y(n20410) );
  NAND2XL U12978 ( .A(n7698), .B(n7697), .Y(n7724) );
  NAND2XL U12979 ( .A(n10426), .B(n10427), .Y(n5003) );
  NAND2X1 U12980 ( .A(n5005), .B(n10425), .Y(n5004) );
  NAND2X1 U12981 ( .A(n10613), .B(n4619), .Y(n10618) );
  NAND2XL U12982 ( .A(n5751), .B(n5298), .Y(n10569) );
  NAND2XL U12983 ( .A(n10564), .B(n10563), .Y(n10592) );
  NOR2XL U12984 ( .A(n15581), .B(n15585), .Y(n15576) );
  NOR2XL U12985 ( .A(n15776), .B(n15775), .Y(n15777) );
  NAND3XL U12986 ( .A(n15826), .B(n15809), .C(n15801), .Y(n15776) );
  NAND4XL U12987 ( .A(n15774), .B(n15827), .C(n15819), .D(n15820), .Y(n15775)
         );
  NOR2XL U12988 ( .A(n15773), .B(n15806), .Y(n15774) );
  NOR4XL U12989 ( .A(n20800), .B(n20791), .C(n23776), .D(n20790), .Y(n9193) );
  XOR2X1 U12990 ( .A(n11797), .B(n5788), .Y(n11821) );
  OAI21XL U12991 ( .A0(n12443), .A1(n12444), .B0(n12442), .Y(n5404) );
  XNOR2X1 U12992 ( .A(n5405), .B(n12443), .Y(n12479) );
  OAI22XL U12993 ( .A0(n12578), .A1(n12577), .B0(n12718), .B1(
        M3_mult_x_15_a_17_), .Y(n12695) );
  INVXL U12994 ( .A(n12807), .Y(n12810) );
  NOR2X1 U12995 ( .A(n14590), .B(n14573), .Y(n14550) );
  XNOR3X2 U12996 ( .A(n5873), .B(n5923), .C(n17590), .Y(n17668) );
  INVXL U12997 ( .A(n18376), .Y(n4870) );
  AOI21XL U12998 ( .A0(n14482), .A1(n14481), .B0(n14480), .Y(n14483) );
  XOR2XL U12999 ( .A(n14479), .B(n14478), .Y(n14481) );
  INVX1 U13000 ( .A(n14663), .Y(n5498) );
  NOR2X1 U13001 ( .A(n14323), .B(n14324), .Y(n14529) );
  INVXL U13002 ( .A(n14529), .Y(n14543) );
  ADDFX2 U13003 ( .A(n12650), .B(n12649), .CI(n12648), .CO(n12680), .S(n12682)
         );
  OR2X2 U13004 ( .A(n12683), .B(n12682), .Y(n5930) );
  NAND2XL U13005 ( .A(n14332), .B(n14331), .Y(n14499) );
  NAND2XL U13006 ( .A(n14535), .B(n14539), .Y(n14487) );
  NOR2X2 U13007 ( .A(n13993), .B(n13992), .Y(n14603) );
  OAI2BB1XL U13008 ( .A0N(n14298), .A1N(n6191), .B0(n23173), .Y(n14304) );
  INVXL U13009 ( .A(n14650), .Y(n14344) );
  NAND2XL U13010 ( .A(n14343), .B(n14342), .Y(n14650) );
  AOI21X1 U13011 ( .A0(n14647), .A1(n14646), .B0(n14645), .Y(n14648) );
  NOR2XL U13012 ( .A(n18721), .B(M3_mult_x_15_b_22_), .Y(n18672) );
  NOR2XL U13013 ( .A(n19960), .B(n19964), .Y(n19955) );
  NAND3XL U13014 ( .A(n25344), .B(n20254), .C(n24828), .Y(n20163) );
  NAND2XL U13015 ( .A(n8756), .B(n8755), .Y(n8757) );
  INVXL U13016 ( .A(n8754), .Y(n8756) );
  NAND2XL U13017 ( .A(n8751), .B(n8750), .Y(n8752) );
  INVXL U13018 ( .A(n8749), .Y(n8751) );
  NAND4XL U13019 ( .A(n9021), .B(n20450), .C(n20449), .D(n20454), .Y(n9022) );
  NOR2XL U13020 ( .A(n9020), .B(n9019), .Y(n9021) );
  NAND3XL U13021 ( .A(n20415), .B(n20432), .C(n20411), .Y(n9020) );
  NAND4XL U13022 ( .A(n9018), .B(n20461), .C(n20435), .D(n20436), .Y(n9019) );
  NAND2XL U13023 ( .A(n20041), .B(n20054), .Y(n20042) );
  INVXL U13024 ( .A(n20055), .Y(n20040) );
  NAND2XL U13025 ( .A(n20044), .B(n20055), .Y(n20045) );
  NOR2XL U13026 ( .A(n15764), .B(n15825), .Y(n15812) );
  INVXL U13027 ( .A(n15820), .Y(n15811) );
  INVXL U13028 ( .A(n15819), .Y(n15822) );
  NAND2XL U13029 ( .A(n21812), .B(n21811), .Y(n22089) );
  INVXL U13030 ( .A(n22085), .Y(n22090) );
  INVXL U13031 ( .A(n22077), .Y(n22092) );
  NOR2XL U13032 ( .A(n23119), .B(n23118), .Y(n21440) );
  NOR2XL U13033 ( .A(n23123), .B(n23122), .Y(n21438) );
  NAND2XL U13034 ( .A(n21176), .B(n21175), .Y(n21790) );
  NAND3XL U13035 ( .A(cs[0]), .B(cs[1]), .C(y20[3]), .Y(n21175) );
  NAND2XL U13036 ( .A(n21355), .B(n21421), .Y(n21358) );
  NAND2XL U13037 ( .A(n21311), .B(temp0[17]), .Y(n21298) );
  NOR2XL U13038 ( .A(n21342), .B(n21520), .Y(n21296) );
  NAND2X1 U13039 ( .A(n21383), .B(n21334), .Y(n21385) );
  AOI21XL U13040 ( .A0(n21207), .A1(n21206), .B0(n21205), .Y(n21234) );
  NOR2XL U13041 ( .A(n21204), .B(n21179), .Y(n21207) );
  NAND2XL U13042 ( .A(n21225), .B(n21469), .Y(n21226) );
  AOI21XL U13043 ( .A0(n21272), .A1(n21271), .B0(n21270), .Y(n21288) );
  NAND2XL U13044 ( .A(n21261), .B(n21473), .Y(n21262) );
  NAND2XL U13045 ( .A(n21279), .B(n21513), .Y(n21280) );
  NOR2XL U13046 ( .A(n21273), .B(n21457), .Y(n21257) );
  NOR2XL U13047 ( .A(n21264), .B(n21245), .Y(n21246) );
  NOR2XL U13048 ( .A(n21470), .B(n21260), .Y(n21245) );
  INVXL U13049 ( .A(n22301), .Y(n22304) );
  NAND2XL U13050 ( .A(n3126), .B(n22302), .Y(n22303) );
  NOR2XL U13051 ( .A(n22203), .B(n22185), .Y(n22135) );
  INVXL U13052 ( .A(n22297), .Y(n22234) );
  NAND2XL U13053 ( .A(n22188), .B(n22301), .Y(n22233) );
  INVXL U13054 ( .A(n22296), .Y(n22299) );
  NAND2XL U13055 ( .A(n3126), .B(n22297), .Y(n22298) );
  INVXL U13056 ( .A(n22295), .Y(n22232) );
  NAND2XL U13057 ( .A(n3126), .B(n22296), .Y(n22231) );
  INVXL U13058 ( .A(n22252), .Y(n22423) );
  AOI21XL U13059 ( .A0(n22295), .A1(n3126), .B0(n22294), .Y(n22344) );
  INVXL U13060 ( .A(n22292), .Y(n22293) );
  AOI2BB1XL U13061 ( .A0N(n22144), .A1N(n22295), .B0(n22292), .Y(n22145) );
  AOI2BB1XL U13062 ( .A0N(n22297), .A1N(n22143), .B0(n22296), .Y(n22144) );
  AOI2BB1XL U13063 ( .A0N(n22142), .A1N(n22302), .B0(n22301), .Y(n22143) );
  AOI2BB1XL U13064 ( .A0N(n22141), .A1N(n22202), .B0(n22305), .Y(n22142) );
  NAND2XL U13065 ( .A(n21918), .B(n21917), .Y(n21919) );
  INVXL U13066 ( .A(n22067), .Y(n22025) );
  AOI21XL U13067 ( .A0(n22048), .A1(n22047), .B0(n22046), .Y(n22049) );
  INVXL U13068 ( .A(n22042), .Y(n22045) );
  NAND2XL U13069 ( .A(n22041), .B(n22047), .Y(n22050) );
  NAND2XL U13070 ( .A(n21965), .B(n21964), .Y(n22053) );
  INVXL U13071 ( .A(n22064), .Y(n22065) );
  NAND2XL U13072 ( .A(n22063), .B(n22066), .Y(n22069) );
  NAND2XL U13073 ( .A(n21927), .B(n21926), .Y(n21928) );
  INVXL U13074 ( .A(n21925), .Y(n21927) );
  NAND2XL U13075 ( .A(n21914), .B(n21913), .Y(n21915) );
  INVXL U13076 ( .A(n21912), .Y(n21914) );
  NAND2XL U13077 ( .A(n21905), .B(n22043), .Y(n21906) );
  INVXL U13078 ( .A(n22044), .Y(n21905) );
  NAND2XL U13079 ( .A(n21935), .B(n21934), .Y(n21936) );
  INVXL U13080 ( .A(n21931), .Y(n21932) );
  INVXL U13081 ( .A(n8977), .Y(n8978) );
  NAND2XL U13082 ( .A(n8976), .B(n8975), .Y(n8980) );
  OAI31XL U13083 ( .A0(n20449), .A1(n20450), .A2(n8974), .B0(n8973), .Y(n8975)
         );
  NAND2XL U13084 ( .A(n14427), .B(y10[24]), .Y(n9118) );
  NAND2XL U13085 ( .A(n14427), .B(y10[26]), .Y(n9125) );
  NAND2XL U13086 ( .A(n14427), .B(y10[30]), .Y(n9110) );
  OAI21XL U13087 ( .A0(n17001), .A1(n17002), .B0(n17000), .Y(n5950) );
  NAND2XL U13088 ( .A(M6_mult_x_15_n483), .B(M6_mult_x_15_n490), .Y(n11358) );
  OR2X2 U13089 ( .A(n7678), .B(n7677), .Y(n7812) );
  NOR2XL U13090 ( .A(n7815), .B(n7746), .Y(n7805) );
  NOR2XL U13091 ( .A(M6_mult_x_15_n582), .B(M6_mult_x_15_n592), .Y(n11109) );
  AOI21XL U13092 ( .A0(n11279), .A1(n11108), .B0(n11107), .Y(n11123) );
  NOR2XL U13093 ( .A(M6_mult_x_15_n593), .B(M6_mult_x_15_n603), .Y(n11119) );
  NAND2XL U13094 ( .A(M6_mult_x_15_n593), .B(M6_mult_x_15_n603), .Y(n11120) );
  NAND2XL U13095 ( .A(M6_mult_x_15_n582), .B(M6_mult_x_15_n592), .Y(n11110) );
  NAND2XL U13096 ( .A(M6_mult_x_15_n482), .B(M6_mult_x_15_n476), .Y(n11350) );
  NOR2XL U13097 ( .A(M6_mult_x_15_n482), .B(M6_mult_x_15_n476), .Y(n10997) );
  NOR2XL U13098 ( .A(n7659), .B(n7658), .Y(n7611) );
  NAND2X1 U13099 ( .A(n20853), .B(n20869), .Y(n20828) );
  NOR2XL U13100 ( .A(M6_mult_x_15_n615), .B(M6_mult_x_15_n625), .Y(n11124) );
  NAND2XL U13101 ( .A(M6_mult_x_15_n615), .B(M6_mult_x_15_n625), .Y(n11276) );
  XOR2X1 U13102 ( .A(n17795), .B(n17797), .Y(n5889) );
  OR2X2 U13103 ( .A(n18590), .B(n18589), .Y(n6093) );
  INVXL U13104 ( .A(n18981), .Y(n18982) );
  INVX1 U13105 ( .A(n17147), .Y(n17146) );
  NOR2X1 U13106 ( .A(n17371), .B(n17144), .Y(n5339) );
  INVX1 U13107 ( .A(n17144), .Y(n5666) );
  NAND2XL U13108 ( .A(n17282), .B(n17281), .Y(n17415) );
  AOI22XL U13109 ( .A0(n17280), .A1(n17279), .B0(n17278), .B1(n18810), .Y(
        n17281) );
  NAND2XL U13110 ( .A(n17283), .B(n17275), .Y(n17282) );
  INVXL U13111 ( .A(n17277), .Y(n17279) );
  NOR2XL U13112 ( .A(n17293), .B(n17292), .Y(n17417) );
  NAND2XL U13113 ( .A(n17291), .B(n17290), .Y(n17292) );
  INVXL U13114 ( .A(n17283), .Y(n17293) );
  XOR2XL U13115 ( .A(n17289), .B(n17288), .Y(n17290) );
  INVXL U13116 ( .A(n20450), .Y(n20419) );
  NAND2XL U13117 ( .A(n3067), .B(n20453), .Y(n20418) );
  XOR2XL U13118 ( .A(n9163), .B(n10671), .Y(n9167) );
  XOR2XL U13119 ( .A(n10676), .B(n10672), .Y(n9156) );
  INVXL U13120 ( .A(n20454), .Y(n20421) );
  NAND2XL U13121 ( .A(n3067), .B(n20457), .Y(n20420) );
  INVXL U13122 ( .A(n9004), .Y(n9008) );
  INVXL U13123 ( .A(n20255), .Y(n20185) );
  OAI21X1 U13124 ( .A0(n10243), .A1(n10242), .B0(n10241), .Y(n10246) );
  NAND2XL U13125 ( .A(n10572), .B(n10571), .Y(n10648) );
  OAI21XL U13126 ( .A0(n10586), .A1(n10591), .B0(n10592), .Y(n10651) );
  INVXL U13127 ( .A(n10666), .Y(n6141) );
  NAND2XL U13128 ( .A(n12796), .B(n12795), .Y(n12830) );
  ADDFX2 U13129 ( .A(n12739), .B(n12738), .CI(n12737), .CO(n12790), .S(n12785)
         );
  INVX1 U13130 ( .A(n12833), .Y(n12853) );
  NOR2X2 U13131 ( .A(n13596), .B(n13595), .Y(n14399) );
  NAND2XL U13132 ( .A(n14383), .B(n14382), .Y(n14480) );
  NAND2XL U13133 ( .A(n14384), .B(n14375), .Y(n14383) );
  AOI22XL U13134 ( .A0(n14381), .A1(n14380), .B0(n14379), .B1(n14378), .Y(
        n14382) );
  XOR2XL U13135 ( .A(n14374), .B(n14373), .Y(n14375) );
  NOR2XL U13136 ( .A(n14396), .B(n14395), .Y(n14482) );
  NAND2BXL U13137 ( .AN(n14394), .B(n14393), .Y(n14395) );
  INVXL U13138 ( .A(n14384), .Y(n14396) );
  XOR2XL U13139 ( .A(n14388), .B(n14387), .Y(n14394) );
  AOI21XL U13140 ( .A0(n18896), .A1(n18865), .B0(n18867), .Y(n18868) );
  NAND4X1 U13141 ( .A(n20321), .B(n13036), .C(n23484), .D(n20317), .Y(n4982)
         );
  NOR4XL U13142 ( .A(n25184), .B(n24087), .C(n24336), .D(n25804), .Y(n11619)
         );
  INVXL U13143 ( .A(n24285), .Y(n11617) );
  NOR2X2 U13144 ( .A(n14639), .B(n14637), .Y(n14629) );
  INVXL U13145 ( .A(n19008), .Y(n19009) );
  INVXL U13146 ( .A(n14514), .Y(n14516) );
  NAND2XL U13147 ( .A(n14511), .B(n14509), .Y(n14507) );
  INVXL U13148 ( .A(temp0[30]), .Y(n7884) );
  NAND2XL U13149 ( .A(n8872), .B(n8871), .Y(n8873) );
  NAND2XL U13150 ( .A(n8866), .B(n8865), .Y(n8867) );
  INVXL U13151 ( .A(n8864), .Y(n8866) );
  NAND2XL U13152 ( .A(n8844), .B(n8843), .Y(n8845) );
  INVXL U13153 ( .A(n8842), .Y(n8844) );
  NAND2XL U13154 ( .A(n8849), .B(n8848), .Y(n8850) );
  INVXL U13155 ( .A(n8847), .Y(n8849) );
  NAND2XL U13156 ( .A(n8878), .B(n8876), .Y(n8840) );
  INVXL U13157 ( .A(n8879), .Y(n8837) );
  NAND2XL U13158 ( .A(n8885), .B(n8884), .Y(n8886) );
  INVXL U13159 ( .A(n8883), .Y(n8885) );
  AOI21XL U13160 ( .A0(n8832), .A1(n8872), .B0(n8831), .Y(n8833) );
  INVXL U13161 ( .A(n8869), .Y(n8832) );
  INVXL U13162 ( .A(n8827), .Y(n8828) );
  INVXL U13163 ( .A(n20254), .Y(n20257) );
  INVXL U13164 ( .A(n24717), .Y(n24678) );
  OAI21XL U13165 ( .A0(n3072), .A1(n20258), .B0(n20240), .Y(n24683) );
  INVXL U13166 ( .A(n24849), .Y(n24826) );
  NOR2XL U13167 ( .A(n24986), .B(n24746), .Y(n24747) );
  INVXL U13168 ( .A(n24798), .Y(n24745) );
  NAND2XL U13169 ( .A(n15730), .B(n15732), .Y(n15703) );
  INVXL U13170 ( .A(n15702), .Y(n15704) );
  AOI31XL U13171 ( .A0(n15721), .A1(n15701), .A2(n15725), .B0(n15700), .Y(
        n15702) );
  INVXL U13172 ( .A(n24871), .Y(n21002) );
  NAND2XL U13173 ( .A(n25269), .B(n21000), .Y(n21001) );
  NAND2XL U13174 ( .A(n15635), .B(n15634), .Y(n15636) );
  INVXL U13175 ( .A(n15633), .Y(n15635) );
  NOR2XL U13176 ( .A(n24916), .B(n24915), .Y(n25011) );
  NOR2XL U13177 ( .A(n15764), .B(n15716), .Y(n24915) );
  INVXL U13178 ( .A(n25270), .Y(n25008) );
  NOR2X1 U13179 ( .A(n22190), .B(n22189), .Y(n22237) );
  NOR2XL U13180 ( .A(n22308), .B(n22141), .Y(n22189) );
  AOI22XL U13181 ( .A0(n21727), .A1(n21718), .B0(n21730), .B1(n21717), .Y(
        n21725) );
  NOR4BXL U13182 ( .AN(n21706), .B(n21705), .C(n21704), .D(n21703), .Y(n21736)
         );
  INVXL U13183 ( .A(n21727), .Y(n21729) );
  INVXL U13184 ( .A(n21730), .Y(n21732) );
  OAI211XL U13185 ( .A0(n21801), .A1(n21682), .B0(n21681), .C0(n21680), .Y(
        n21695) );
  NOR2XL U13186 ( .A(n21685), .B(n21684), .Y(n21686) );
  AOI21XL U13187 ( .A0(n21687), .A1(n21507), .B0(n21683), .Y(n21685) );
  NAND2XL U13188 ( .A(n21331), .B(w1[26]), .Y(n21323) );
  AOI211XL U13189 ( .A0(n15725), .A1(n15724), .B0(n15872), .C0(n15873), .Y(
        n15727) );
  AOI211XL U13190 ( .A0(n15720), .A1(n15719), .B0(n15819), .C0(n15820), .Y(
        n15723) );
  NAND2XL U13191 ( .A(n15474), .B(n15473), .Y(n15475) );
  INVXL U13192 ( .A(n15472), .Y(n15474) );
  NAND2XL U13193 ( .A(n15465), .B(n15605), .Y(n15466) );
  INVXL U13194 ( .A(n15606), .Y(n15465) );
  NOR2XL U13195 ( .A(n22308), .B(n22277), .Y(n22278) );
  NOR2XL U13196 ( .A(n22249), .B(n22248), .Y(n22324) );
  NOR2XL U13197 ( .A(n22308), .B(n22276), .Y(n22248) );
  INVXL U13198 ( .A(n22273), .Y(n22246) );
  AOI22XL U13199 ( .A0(n22344), .A1(n22343), .B0(n22342), .B1(n3129), .Y(
        n22351) );
  NAND2XL U13200 ( .A(n22060), .B(n22059), .Y(n22061) );
  NAND2XL U13201 ( .A(n21333), .B(w1[24]), .Y(n21303) );
  NAND2XL U13202 ( .A(n21331), .B(w1[28]), .Y(n21316) );
  INVXL U13203 ( .A(n22015), .Y(n22016) );
  INVXL U13204 ( .A(n22057), .Y(n22020) );
  NAND2XL U13205 ( .A(n19346), .B(w2[24]), .Y(n8076) );
  NAND3BXL U13206 ( .AN(n11100), .B(n20725), .C(n20291), .Y(n11382) );
  NAND4XL U13207 ( .A(n20625), .B(n23916), .C(n20290), .D(n11465), .Y(n11100)
         );
  NAND2XL U13208 ( .A(n23498), .B(n23896), .Y(n11383) );
  NAND3BXL U13209 ( .AN(n9186), .B(n23661), .C(n24383), .Y(n9187) );
  NAND4XL U13210 ( .A(n24269), .B(n20800), .C(n20791), .D(n23776), .Y(n9186)
         );
  NAND2XL U13211 ( .A(n14427), .B(y10[27]), .Y(n9130) );
  NAND2XL U13212 ( .A(n25233), .B(sigma10[27]), .Y(n9131) );
  NAND2XL U13213 ( .A(n4826), .B(y12[27]), .Y(n9129) );
  NAND2XL U13214 ( .A(n14427), .B(y10[23]), .Y(n9114) );
  NAND2XL U13215 ( .A(n4856), .B(target_temp[29]), .Y(n14432) );
  NOR2XL U13216 ( .A(n23503), .B(n23501), .Y(n23497) );
  XOR2XL U13217 ( .A(n10996), .B(n10995), .Y(n23498) );
  NAND2XL U13218 ( .A(n10994), .B(n10993), .Y(n10995) );
  AOI21XL U13219 ( .A0(n11099), .A1(n11097), .B0(n10991), .Y(n10996) );
  INVXL U13220 ( .A(n10992), .Y(n10994) );
  NAND2XL U13221 ( .A(n23896), .B(n23895), .Y(n20769) );
  XNOR2XL U13222 ( .A(n10977), .B(n10976), .Y(n20766) );
  NAND2XL U13223 ( .A(n10975), .B(n10974), .Y(n10976) );
  INVXL U13224 ( .A(n10973), .Y(n10975) );
  NAND2XL U13225 ( .A(n7832), .B(n7831), .Y(n7833) );
  INVXL U13226 ( .A(n17391), .Y(n17393) );
  INVXL U13227 ( .A(n17361), .Y(n17363) );
  INVX1 U13228 ( .A(n17326), .Y(n17344) );
  AOI21XL U13229 ( .A0(n11368), .A1(n11367), .B0(n11366), .Y(n11369) );
  INVXL U13230 ( .A(n11365), .Y(n11366) );
  INVXL U13231 ( .A(n11364), .Y(n11368) );
  NOR2XL U13232 ( .A(n19081), .B(n19063), .Y(n23467) );
  XNOR2XL U13233 ( .A(n11105), .B(n11104), .Y(n23468) );
  NAND2XL U13234 ( .A(n11103), .B(n11102), .Y(n11104) );
  INVXL U13235 ( .A(n11101), .Y(n11103) );
  INVX1 U13236 ( .A(n17206), .Y(n6144) );
  INVXL U13237 ( .A(M4_U3_U1_enc_tree_0__4__16_), .Y(n18839) );
  INVXL U13238 ( .A(M4_U3_U1_enc_tree_0__2__12_), .Y(
        M4_U3_U1_enc_tree_0__3__8_) );
  INVXL U13239 ( .A(M4_U4_U1_enc_tree_0__2__12_), .Y(
        M3_U4_U1_enc_tree_0__3__8_) );
  OR2XL U13240 ( .A(M3_U4_U1_or2_tree_0__2__16_), .B(
        M3_U4_U1_or2_tree_0__2__24_), .Y(n26157) );
  NAND2XL U13241 ( .A(n18815), .B(n18814), .Y(n18841) );
  AOI22XL U13242 ( .A0(n18813), .A1(n18812), .B0(n18811), .B1(n18810), .Y(
        n18814) );
  NAND2XL U13243 ( .A(n18816), .B(n18807), .Y(n18815) );
  INVXL U13244 ( .A(n18809), .Y(n18812) );
  NOR2XL U13245 ( .A(n18828), .B(n18827), .Y(n18843) );
  NAND2XL U13246 ( .A(n18826), .B(n18825), .Y(n18827) );
  INVXL U13247 ( .A(n18816), .Y(n18828) );
  XOR2XL U13248 ( .A(n18824), .B(n18823), .Y(n18825) );
  NAND2XL U13249 ( .A(n11011), .B(n11009), .Y(n10957) );
  INVXL U13250 ( .A(n11363), .Y(n11026) );
  INVXL U13251 ( .A(n11371), .Y(n11025) );
  NAND2XL U13252 ( .A(n11412), .B(n23674), .Y(n11447) );
  NAND2XL U13253 ( .A(n23668), .B(n11407), .Y(n11448) );
  AOI21XL U13254 ( .A0(n23678), .A1(n23677), .B0(n6218), .Y(n11407) );
  NAND2XL U13255 ( .A(n21166), .B(sigma10[26]), .Y(n11564) );
  AOI2BB1XL U13256 ( .A0N(n20553), .A1N(n20473), .B0(n20597), .Y(n20554) );
  NAND2XL U13257 ( .A(n7818), .B(n7816), .Y(n7803) );
  AOI21XL U13258 ( .A0(n9181), .A1(n9160), .B0(n9162), .Y(n9174) );
  INVXL U13259 ( .A(n9179), .Y(n9162) );
  NOR2XL U13260 ( .A(n9167), .B(n10694), .Y(n9170) );
  NAND2XL U13261 ( .A(n9167), .B(n10694), .Y(n9171) );
  NOR2XL U13262 ( .A(n10693), .B(n9156), .Y(n9175) );
  NAND2XL U13263 ( .A(n10693), .B(n9156), .Y(n9176) );
  AOI2BB2XL U13264 ( .B0(n20499), .B1(n20473), .A0N(n20535), .A1N(n20473), .Y(
        n20598) );
  NAND2XL U13265 ( .A(n9133), .B(n14413), .Y(n9134) );
  NAND2XL U13266 ( .A(n25233), .B(sigma10[28]), .Y(n9133) );
  INVX1 U13267 ( .A(n19315), .Y(n19294) );
  INVXL U13268 ( .A(n19333), .Y(n19336) );
  INVXL U13269 ( .A(n19329), .Y(n19332) );
  OAI21X1 U13270 ( .A0(n19564), .A1(n19328), .B0(n19327), .Y(n23210) );
  INVXL U13271 ( .A(n19325), .Y(n19328) );
  OAI21XL U13272 ( .A0(n3068), .A1(n20508), .B0(n20507), .Y(n20524) );
  OAI21XL U13273 ( .A0(n20473), .A1(n20494), .B0(n20478), .Y(n20517) );
  NOR2XL U13274 ( .A(n20583), .B(n3071), .Y(n20584) );
  NOR2XL U13275 ( .A(n20582), .B(n20581), .Y(n20585) );
  NOR2XL U13276 ( .A(n3124), .B(n20580), .Y(n20581) );
  NOR2XL U13277 ( .A(n3067), .B(n20579), .Y(n20582) );
  INVX1 U13278 ( .A(n19334), .Y(n19301) );
  INVXL U13279 ( .A(n14938), .Y(n14941) );
  NAND2XL U13280 ( .A(n7718), .B(n7723), .Y(n7719) );
  INVXL U13281 ( .A(n7725), .Y(n7718) );
  INVXL U13282 ( .A(n10623), .Y(n10625) );
  OAI21X1 U13283 ( .A0(n5237), .A1(n10647), .B0(n10636), .Y(n4859) );
  INVXL U13284 ( .A(n10582), .Y(n10584) );
  INVXL U13285 ( .A(n20614), .Y(n20703) );
  OAI21XL U13286 ( .A0(n12846), .A1(n12848), .B0(n12849), .Y(n5400) );
  OAI21XL U13287 ( .A0(n26297), .A1(n3115), .B0(n14411), .Y(n14697) );
  NAND2XL U13288 ( .A(in_valid_t), .B(w2[59]), .Y(n18750) );
  NAND2XL U13289 ( .A(n3111), .B(data[91]), .Y(n18752) );
  INVXL U13290 ( .A(n20653), .Y(n6147) );
  INVX1 U13291 ( .A(n19311), .Y(n19296) );
  INVXL U13292 ( .A(temp0[23]), .Y(n8066) );
  INVX1 U13293 ( .A(n8189), .Y(n8163) );
  AOI2BB2XL U13294 ( .B0(n20259), .B1(n3069), .A0N(n20231), .A1N(n3069), .Y(
        n24752) );
  NAND2XL U13295 ( .A(n20115), .B(n20117), .Y(n20081) );
  INVXL U13296 ( .A(n20080), .Y(n20082) );
  AOI31XL U13297 ( .A0(n20106), .A1(n20079), .A2(n20110), .B0(n20078), .Y(
        n20080) );
  AOI2BB2XL U13298 ( .B0(n20259), .B1(n20182), .A0N(n24751), .A1N(n20182), .Y(
        n24898) );
  NAND2XL U13299 ( .A(n24895), .B(n24894), .Y(n24896) );
  AOI2BB2XL U13300 ( .B0(n24825), .B1(n3069), .A0N(n24683), .A1N(n3069), .Y(
        n24994) );
  NOR2XL U13301 ( .A(n24988), .B(n24987), .Y(n24991) );
  NOR2XL U13302 ( .A(n24989), .B(n3032), .Y(n24990) );
  NOR2XL U13303 ( .A(n24986), .B(n20100), .Y(n24987) );
  NAND2XL U13304 ( .A(n3075), .B(n24684), .Y(n24998) );
  NAND2X1 U13305 ( .A(n15849), .B(n3077), .Y(n15916) );
  NAND2XL U13306 ( .A(n21329), .B(temp0[25]), .Y(n21322) );
  OAI21XL U13307 ( .A0(n26145), .A1(n21333), .B0(n21324), .Y(n21434) );
  NAND2XL U13308 ( .A(n21333), .B(temp0[26]), .Y(n21324) );
  OAI21X1 U13309 ( .A0(n21519), .A1(n21424), .B0(n21423), .Y(n23125) );
  INVXL U13310 ( .A(n21421), .Y(n21424) );
  NAND2XL U13311 ( .A(n21393), .B(n21422), .Y(n21423) );
  NAND2XL U13312 ( .A(n23282), .B(n23277), .Y(n22407) );
  OAI21XL U13313 ( .A0(n6170), .A1(n21333), .B0(n21317), .Y(n21409) );
  NAND2XL U13314 ( .A(n21331), .B(temp0[28]), .Y(n21317) );
  NOR3X1 U13315 ( .A(n23412), .B(n23393), .C(n22176), .Y(n22173) );
  INVXL U13316 ( .A(n22258), .Y(n22215) );
  INVXL U13317 ( .A(n22213), .Y(n22214) );
  INVXL U13318 ( .A(n19034), .Y(n19036) );
  NOR2XL U13319 ( .A(n19030), .B(n19029), .Y(n19039) );
  INVXL U13320 ( .A(n19028), .Y(n19030) );
  NOR2XL U13321 ( .A(n19033), .B(n19032), .Y(n19038) );
  INVXL U13322 ( .A(n19031), .Y(n19033) );
  NAND2XL U13323 ( .A(n10695), .B(n9161), .Y(n9179) );
  INVXL U13324 ( .A(n10686), .Y(n10689) );
  NAND3XL U13325 ( .A(n10698), .B(n10697), .C(n10696), .Y(n10699) );
  INVXL U13326 ( .A(n10694), .Y(n10697) );
  INVXL U13327 ( .A(n10695), .Y(n10696) );
  NOR2XL U13328 ( .A(n10693), .B(n10692), .Y(n10698) );
  NAND2XL U13329 ( .A(n3223), .B(learning_rate[26]), .Y(n9166) );
  AOI22XL U13330 ( .A0(n25233), .A1(data[26]), .B0(in_valid_d), .B1(w1[282]), 
        .Y(n9165) );
  AOI22XL U13331 ( .A0(n25233), .A1(data[27]), .B0(in_valid_d), .B1(w1[283]), 
        .Y(n9150) );
  NAND2XL U13332 ( .A(n3223), .B(learning_rate[28]), .Y(n9148) );
  AOI22XL U13333 ( .A0(n25233), .A1(data[28]), .B0(in_valid_d), .B1(w1[284]), 
        .Y(n9147) );
  NOR2XL U13334 ( .A(n17401), .B(n17400), .Y(n17410) );
  INVXL U13335 ( .A(n17399), .Y(n17401) );
  NAND2X1 U13336 ( .A(n5100), .B(n20761), .Y(n20764) );
  XOR2XL U13337 ( .A(n23543), .B(n23542), .Y(n23939) );
  INVXL U13338 ( .A(n23541), .Y(n23542) );
  NAND2XL U13339 ( .A(n23915), .B(n23540), .Y(n23543) );
  XOR2X1 U13340 ( .A(n10743), .B(n20275), .Y(n23620) );
  NAND2X1 U13341 ( .A(n5100), .B(n20831), .Y(n20833) );
  INVXL U13342 ( .A(n17450), .Y(n20341) );
  XOR2XL U13343 ( .A(n11584), .B(n13009), .Y(n11614) );
  NAND2XL U13344 ( .A(n24047), .B(n24046), .Y(n24049) );
  INVXL U13345 ( .A(n24045), .Y(n24047) );
  NOR2XL U13346 ( .A(n23802), .B(n23799), .Y(n20603) );
  OAI21XL U13347 ( .A0(n20519), .A1(n3073), .B0(n20424), .Y(n20608) );
  NAND2XL U13348 ( .A(n20423), .B(n20422), .Y(n20424) );
  NAND2XL U13349 ( .A(n20426), .B(n20597), .Y(n20422) );
  NAND2XL U13350 ( .A(in_valid_t), .B(learning_rate[24]), .Y(n11597) );
  NAND2XL U13351 ( .A(n25206), .B(sigma10[24]), .Y(n11599) );
  NAND2XL U13352 ( .A(n19564), .B(n19318), .Y(n19291) );
  AOI2BB2XL U13353 ( .B0(n3030), .B1(n24310), .A0N(n24310), .A1N(n20125), .Y(
        n24308) );
  NAND2X1 U13354 ( .A(n5600), .B(n5100), .Y(n20285) );
  XOR2XL U13355 ( .A(n7397), .B(n7841), .Y(n7407) );
  INVXL U13356 ( .A(n20996), .Y(n24527) );
  NOR2XL U13357 ( .A(n24998), .B(n23200), .Y(n24531) );
  INVX1 U13358 ( .A(n23739), .Y(n5749) );
  INVX1 U13359 ( .A(n17484), .Y(n10716) );
  NAND2X1 U13360 ( .A(n3132), .B(n10715), .Y(n10717) );
  NAND2X1 U13361 ( .A(n3132), .B(n23532), .Y(n5767) );
  INVXL U13362 ( .A(n17485), .Y(n19047) );
  OAI22XL U13363 ( .A0(n25280), .A1(n3076), .B0(n25279), .B1(n25278), .Y(
        n25291) );
  NOR2XL U13364 ( .A(n25277), .B(n25276), .Y(n25278) );
  NOR2XL U13365 ( .A(n25265), .B(n3077), .Y(n25279) );
  AOI2BB2XL U13366 ( .B0(n25269), .B1(n23965), .A0N(n23965), .A1N(n25269), .Y(
        n23964) );
  NAND2X1 U13367 ( .A(n3132), .B(n19073), .Y(n5483) );
  INVXL U13368 ( .A(n12909), .Y(n12911) );
  NAND2X1 U13369 ( .A(n23744), .B(n20329), .Y(n20332) );
  NOR2XL U13370 ( .A(n4294), .B(n20328), .Y(n20329) );
  NAND2XL U13371 ( .A(n23744), .B(n20304), .Y(n20306) );
  NOR2X1 U13372 ( .A(n23709), .B(n20661), .Y(n20662) );
  CLKINVX3 U13373 ( .A(n13026), .Y(n23651) );
  INVXL U13374 ( .A(n23445), .Y(n20974) );
  NOR2XL U13375 ( .A(n23445), .B(n23444), .Y(n23446) );
  XOR2X2 U13376 ( .A(n20665), .B(n5027), .Y(n23702) );
  AND2X2 U13377 ( .A(n23744), .B(n20303), .Y(n5027) );
  NAND3X1 U13378 ( .A(n3357), .B(n5764), .C(n5644), .Y(n5643) );
  NOR2BX1 U13379 ( .AN(n20920), .B(n3958), .Y(n5644) );
  NOR2X1 U13380 ( .A(n20929), .B(n20923), .Y(n5764) );
  OAI21X2 U13381 ( .A0(n19014), .A1(n18958), .B0(n18957), .Y(n5890) );
  NAND2X1 U13382 ( .A(n23744), .B(n23588), .Y(n23591) );
  NAND2X1 U13383 ( .A(n23734), .B(n23457), .Y(n5920) );
  NOR2XL U13384 ( .A(n23478), .B(n23476), .Y(n23457) );
  CMPR32X1 U13385 ( .A(n14711), .B(n14464), .C(n14463), .CO(n14459), .S(n24331) );
  XOR2XL U13386 ( .A(n18763), .B(n19034), .Y(n18772) );
  XOR2XL U13387 ( .A(n14437), .B(n14704), .Y(n14466) );
  AOI2BB2XL U13388 ( .B0(n3067), .B1(n23761), .A0N(n23761), .A1N(n3067), .Y(
        n23759) );
  NOR2XL U13389 ( .A(n20246), .B(n3075), .Y(n20247) );
  AOI21XL U13390 ( .A0(n20066), .A1(n20243), .B0(n20242), .Y(n24611) );
  NOR2XL U13391 ( .A(n24833), .B(n20066), .Y(n20242) );
  NOR2XL U13392 ( .A(n20252), .B(n3075), .Y(n20253) );
  INVXL U13393 ( .A(n24630), .Y(n24645) );
  OAI22XL U13394 ( .A0(n25352), .A1(n3074), .B0(n25351), .B1(n25350), .Y(
        n25362) );
  NOR2XL U13395 ( .A(n25349), .B(n25348), .Y(n25350) );
  AND2XL U13396 ( .A(n25356), .B(n25355), .Y(n25357) );
  NOR2XL U13397 ( .A(n15899), .B(n3077), .Y(n15870) );
  NAND2XL U13398 ( .A(n3079), .B(n22403), .Y(n22399) );
  NOR2XL U13399 ( .A(n22396), .B(n22395), .Y(n22401) );
  NAND2XL U13400 ( .A(n22404), .B(n22403), .Y(n22405) );
  INVXL U13401 ( .A(n23270), .Y(n23268) );
  NAND2XL U13402 ( .A(n23275), .B(n23272), .Y(n23267) );
  NOR2XL U13403 ( .A(n22435), .B(n23113), .Y(n23290) );
  NOR2XL U13404 ( .A(n22385), .B(n22124), .Y(n22388) );
  NOR2XL U13405 ( .A(n23238), .B(n23293), .Y(n23240) );
  NAND2XL U13406 ( .A(n23236), .B(n23265), .Y(n23238) );
  INVXL U13407 ( .A(n23261), .Y(n23236) );
  NAND2X1 U13408 ( .A(n23228), .B(n22216), .Y(n22228) );
  NOR2XL U13409 ( .A(n3079), .B(n3082), .Y(n23114) );
  NOR2XL U13410 ( .A(n22462), .B(n23113), .Y(n23282) );
  NAND2XL U13411 ( .A(n23278), .B(n23277), .Y(n23280) );
  NOR2XL U13412 ( .A(n22380), .B(n23113), .Y(n23285) );
  INVXL U13413 ( .A(n23285), .Y(n23292) );
  NAND2XL U13414 ( .A(n22382), .B(n22461), .Y(n22383) );
  NOR2XL U13415 ( .A(n23293), .B(n23292), .Y(n23295) );
  NOR2XL U13416 ( .A(n23293), .B(n23261), .Y(n23263) );
  NOR2XL U13417 ( .A(n22410), .B(n3082), .Y(n22369) );
  NOR2XL U13418 ( .A(n22433), .B(n22124), .Y(n22376) );
  NOR2XL U13419 ( .A(n22393), .B(n3082), .Y(n22366) );
  NOR2XL U13420 ( .A(n22444), .B(n22124), .Y(n22365) );
  INVXL U13421 ( .A(n23316), .Y(n23343) );
  INVXL U13422 ( .A(n23344), .Y(n23313) );
  NOR2XL U13423 ( .A(n22447), .B(n22124), .Y(n22358) );
  NAND2XL U13424 ( .A(n23346), .B(n23345), .Y(n23348) );
  NOR2XL U13425 ( .A(n23344), .B(n23343), .Y(n23345) );
  INVXL U13426 ( .A(n23341), .Y(n23338) );
  NAND2XL U13427 ( .A(n23307), .B(n23346), .Y(n23309) );
  NOR2XL U13428 ( .A(n23330), .B(n23338), .Y(n23307) );
  OAI22X1 U13429 ( .A0(n22330), .A1(n22329), .B0(n22389), .B1(n22418), .Y(
        n23335) );
  NOR2XL U13430 ( .A(n22328), .B(n22327), .Y(n22329) );
  NAND2XL U13431 ( .A(n23331), .B(n23346), .Y(n23333) );
  INVXL U13432 ( .A(n22386), .Y(n22349) );
  NAND2XL U13433 ( .A(n22347), .B(n22346), .Y(n22348) );
  NAND2XL U13434 ( .A(n23301), .B(n23346), .Y(n23303) );
  NOR2XL U13435 ( .A(n23330), .B(n23300), .Y(n23301) );
  NAND2XL U13436 ( .A(n23299), .B(n23335), .Y(n23300) );
  INVXL U13437 ( .A(n23329), .Y(n23299) );
  INVXL U13438 ( .A(n22410), .Y(n22419) );
  NAND2XL U13439 ( .A(n22416), .B(n22415), .Y(n22417) );
  NAND2XL U13440 ( .A(n22431), .B(n22430), .Y(n22432) );
  OR2XL U13441 ( .A(n22442), .B(n22441), .Y(n22443) );
  INVXL U13442 ( .A(n23369), .Y(n23370) );
  NAND2XL U13443 ( .A(n23383), .B(n23382), .Y(n23385) );
  NAND2XL U13444 ( .A(n21166), .B(target_temp[27]), .Y(n11586) );
  NAND2XL U13445 ( .A(n4875), .B(sigma10[27]), .Y(n11587) );
  NAND2XL U13446 ( .A(n5015), .B(data[123]), .Y(n17172) );
  NAND2X1 U13447 ( .A(in_valid_t), .B(learning_rate[30]), .Y(n11549) );
  INVXL U13448 ( .A(temp0[25]), .Y(n23789) );
  NAND4XL U13449 ( .A(n7857), .B(n7856), .C(n7859), .D(n7858), .Y(n7837) );
  NAND4XL U13450 ( .A(n7853), .B(n7852), .C(n7855), .D(n7854), .Y(n7838) );
  NAND4XL U13451 ( .A(n7863), .B(n7862), .C(n7861), .D(n7860), .Y(n7864) );
  NAND3XL U13452 ( .A(n7851), .B(n7850), .C(n7849), .Y(n7865) );
  NAND4XL U13453 ( .A(n14716), .B(n14710), .C(n14709), .D(n14715), .Y(n14696)
         );
  NAND4XL U13454 ( .A(n14712), .B(n14711), .C(n14714), .D(n14713), .Y(n14695)
         );
  NAND2XL U13455 ( .A(n14693), .B(n14703), .Y(n14694) );
  NAND4XL U13456 ( .A(n17411), .B(n17410), .C(n17409), .D(n17408), .Y(n17412)
         );
  NOR2XL U13457 ( .A(n17404), .B(n17403), .Y(n17409) );
  NOR2XL U13458 ( .A(n17407), .B(n17406), .Y(n17408) );
  NOR2XL U13459 ( .A(n23920), .B(n3115), .Y(n23922) );
  NOR2XL U13460 ( .A(n23505), .B(n3115), .Y(n23507) );
  AOI22XL U13461 ( .A0(n23949), .A1(n23946), .B0(n23947), .B1(n23928), .Y(
        n23505) );
  NOR2XL U13462 ( .A(n23950), .B(n3115), .Y(n23952) );
  AOI22XL U13463 ( .A0(n23949), .A1(n23948), .B0(n23947), .B1(n23946), .Y(
        n23950) );
  AND2X2 U13464 ( .A(n17422), .B(n3357), .Y(n5708) );
  NOR2XL U13465 ( .A(n20300), .B(n3115), .Y(n20301) );
  NOR2XL U13466 ( .A(n23929), .B(n3115), .Y(n23930) );
  NOR2XL U13467 ( .A(n23727), .B(n3115), .Y(n23729) );
  NOR2XL U13468 ( .A(n23934), .B(n3115), .Y(n23936) );
  NOR2XL U13469 ( .A(n23908), .B(n3115), .Y(n23910) );
  NOR2XL U13470 ( .A(n20773), .B(n3115), .Y(n20774) );
  NOR2XL U13471 ( .A(n23887), .B(n9146), .Y(n23889) );
  NOR2XL U13472 ( .A(n20825), .B(n9146), .Y(n20826) );
  NAND3X1 U13473 ( .A(n19104), .B(n23521), .C(in_valid_d), .Y(n5205) );
  NAND3X1 U13474 ( .A(n23522), .B(n3128), .C(in_valid_d), .Y(n5206) );
  NOR2XL U13475 ( .A(n19084), .B(n3115), .Y(n19086) );
  NOR2XL U13476 ( .A(n23900), .B(n9146), .Y(n23901) );
  NOR2XL U13477 ( .A(n20963), .B(n9146), .Y(n20964) );
  OR2XL U13478 ( .A(n20958), .B(n20957), .Y(n20960) );
  NAND3BX1 U13479 ( .AN(n17468), .B(n4653), .C(n3357), .Y(n5709) );
  NAND2X1 U13480 ( .A(n4653), .B(n5393), .Y(n5696) );
  NOR2XL U13481 ( .A(n5697), .B(n17468), .Y(n5393) );
  NOR2X1 U13482 ( .A(n20929), .B(n20355), .Y(n20356) );
  NOR2X1 U13483 ( .A(n20929), .B(n20358), .Y(n20359) );
  XOR2XL U13484 ( .A(n20723), .B(n20722), .Y(n20730) );
  INVXL U13485 ( .A(n20721), .Y(n20722) );
  NAND2XL U13486 ( .A(n23915), .B(n20720), .Y(n20723) );
  NAND2XL U13487 ( .A(n5874), .B(n6091), .Y(n4643) );
  NOR2XL U13488 ( .A(n20628), .B(n3115), .Y(n20630) );
  AOI22XL U13489 ( .A0(n25725), .A1(n23949), .B0(n23947), .B1(n20627), .Y(
        n20628) );
  NOR2XL U13490 ( .A(n20728), .B(n3115), .Y(n25724) );
  XOR2XL U13491 ( .A(n20727), .B(n20726), .Y(n25727) );
  INVXL U13492 ( .A(n20725), .Y(n20726) );
  NAND2XL U13493 ( .A(n23915), .B(n20724), .Y(n20727) );
  NOR2XL U13494 ( .A(n20717), .B(n3115), .Y(n25728) );
  XOR2X1 U13495 ( .A(n17438), .B(n4855), .Y(n17448) );
  OAI2BB1XL U13496 ( .A0N(n25701), .A1N(n25700), .B0(n25699), .Y(n25702) );
  INVXL U13497 ( .A(n23608), .Y(n23605) );
  AOI22X1 U13498 ( .A0(n20385), .A1(n4779), .B0(n24792), .B1(n25300), .Y(
        n25319) );
  INVXL U13499 ( .A(n24769), .Y(n20776) );
  INVX2 U13500 ( .A(n3455), .Y(n5586) );
  NOR2X1 U13501 ( .A(n20804), .B(n20803), .Y(n25842) );
  INVXL U13502 ( .A(n23661), .Y(n20798) );
  INVX1 U13503 ( .A(n24386), .Y(n5229) );
  NOR2X1 U13504 ( .A(n24388), .B(n24387), .Y(n24449) );
  INVXL U13505 ( .A(n24383), .Y(n24381) );
  NOR2X1 U13506 ( .A(n24273), .B(n24272), .Y(n25093) );
  INVXL U13507 ( .A(n24270), .Y(n24271) );
  NAND2XL U13508 ( .A(n23255), .B(n22464), .Y(n23038) );
  AOI22XL U13509 ( .A0(n3100), .A1(n23202), .B0(n3041), .B1(n23201), .Y(n23215) );
  AOI2BB1XL U13510 ( .A0N(n24067), .A1N(n23213), .B0(n3215), .Y(n23214) );
  INVXL U13511 ( .A(n24065), .Y(n23216) );
  AOI22X1 U13512 ( .A0(n20385), .A1(n20877), .B0(n25300), .B1(n20876), .Y(
        n23656) );
  INVXL U13513 ( .A(n20877), .Y(n20874) );
  AOI22X1 U13514 ( .A0(n20385), .A1(n20906), .B0(n25300), .B1(n20905), .Y(
        n24642) );
  INVXL U13515 ( .A(n23754), .Y(n23752) );
  AOI22X1 U13516 ( .A0(n20385), .A1(n24712), .B0(n24711), .B1(n25300), .Y(
        n25316) );
  INVXL U13517 ( .A(n24712), .Y(n24709) );
  INVX1 U13518 ( .A(n20914), .Y(n24490) );
  OAI2BB1X1 U13519 ( .A0N(n23868), .A1N(n23867), .B0(n23866), .Y(n25707) );
  OAI2BB1X1 U13520 ( .A0N(n23868), .A1N(n23824), .B0(n23823), .Y(n25720) );
  AOI21XL U13521 ( .A0(n23864), .A1(n23822), .B0(n23863), .Y(n23823) );
  AOI22X2 U13522 ( .A0(n23741), .A1(n3128), .B0(n23945), .B1(n19104), .Y(
        n24656) );
  INVXL U13523 ( .A(n24860), .Y(n24815) );
  AOI22X2 U13524 ( .A0(n20716), .A1(n19104), .B0(n5523), .B1(n3128), .Y(n25747) );
  CLKINVX3 U13525 ( .A(n24380), .Y(n5353) );
  INVXL U13526 ( .A(n20946), .Y(n20948) );
  NOR2XL U13527 ( .A(n20945), .B(n20944), .Y(n20946) );
  NAND2XL U13528 ( .A(n5269), .B(n24206), .Y(n5821) );
  NAND2X1 U13529 ( .A(n24210), .B(n24117), .Y(n5879) );
  AOI22X1 U13530 ( .A0(n3081), .A1(n23793), .B0(n23792), .B1(n4267), .Y(n24715) );
  NAND2X1 U13531 ( .A(n23792), .B(n23883), .Y(n5271) );
  AOI22X2 U13532 ( .A0(n23702), .A1(n4267), .B0(n3081), .B1(n23703), .Y(n24796) );
  INVXL U13533 ( .A(n24160), .Y(n4966) );
  NAND2X1 U13534 ( .A(n25378), .B(n5428), .Y(n5427) );
  INVX1 U13535 ( .A(n24256), .Y(n5428) );
  NOR2X1 U13536 ( .A(n3014), .B(n23550), .Y(n5772) );
  NAND2X2 U13537 ( .A(n5911), .B(n24111), .Y(n6022) );
  AOI21X1 U13538 ( .A0(n5911), .A1(n25126), .B0(n5866), .Y(n25783) );
  XOR2XL U13539 ( .A(n25125), .B(n25129), .Y(n25126) );
  NAND2X1 U13540 ( .A(n6085), .B(n6132), .Y(n5866) );
  NAND2X1 U13541 ( .A(n25128), .B(n25129), .Y(n6085) );
  INVXL U13542 ( .A(n23809), .Y(n23813) );
  INVXL U13543 ( .A(n23815), .Y(n23819) );
  INVXL U13544 ( .A(n23689), .Y(n23693) );
  INVX1 U13545 ( .A(n23836), .Y(n25393) );
  INVX1 U13546 ( .A(n25030), .Y(n25372) );
  INVXL U13547 ( .A(n23869), .Y(n23875) );
  INVXL U13548 ( .A(n9029), .Y(n9037) );
  INVX1 U13549 ( .A(n24612), .Y(n25518) );
  AOI22XL U13550 ( .A0(n24692), .A1(n24611), .B0(n24908), .B1(n24610), .Y(
        n24612) );
  INVXL U13551 ( .A(n24611), .Y(n24608) );
  INVX1 U13552 ( .A(n24463), .Y(n25677) );
  AOI22XL U13553 ( .A0(n24692), .A1(n24462), .B0(n24908), .B1(n24461), .Y(
        n24463) );
  AOI22XL U13554 ( .A0(n24692), .A1(n20683), .B0(n24908), .B1(n20682), .Y(
        n20684) );
  AOI22XL U13555 ( .A0(n24692), .A1(n24492), .B0(n24908), .B1(n24478), .Y(
        n24479) );
  INVXL U13556 ( .A(n24492), .Y(n24477) );
  INVX1 U13557 ( .A(n24693), .Y(n25472) );
  AOI22XL U13558 ( .A0(n24692), .A1(n24726), .B0(n24908), .B1(n24691), .Y(
        n24693) );
  XOR2XL U13559 ( .A(n24690), .B(n24687), .Y(n24691) );
  INVXL U13560 ( .A(n24807), .Y(n24762) );
  AOI22XL U13561 ( .A0(n24692), .A1(n24859), .B0(n24908), .B1(n24838), .Y(
        n24839) );
  INVXL U13562 ( .A(n24859), .Y(n24836) );
  NAND2XL U13563 ( .A(n24503), .B(n24502), .Y(n24505) );
  INVXL U13564 ( .A(n24584), .Y(n24556) );
  INVXL U13565 ( .A(n24591), .Y(n24588) );
  NOR2XL U13566 ( .A(n24587), .B(n24586), .Y(n24589) );
  INVXL U13567 ( .A(n24618), .Y(n24602) );
  INVXL U13568 ( .A(n24771), .Y(n15904) );
  INVXL U13569 ( .A(n24780), .Y(n24777) );
  AOI22XL U13570 ( .A0(n3029), .A1(n24975), .B0(n25290), .B1(n24884), .Y(
        n25408) );
  INVXL U13571 ( .A(n24977), .Y(n24882) );
  INVXL U13572 ( .A(n24974), .Y(n24930) );
  NAND2X1 U13573 ( .A(in_valid_d), .B(data_point[23]), .Y(n24022) );
  NAND2X1 U13574 ( .A(in_valid_d), .B(data_point[25]), .Y(n25216) );
  NAND2X1 U13575 ( .A(in_valid_d), .B(data_point[27]), .Y(n25213) );
  NAND2X1 U13576 ( .A(in_valid_d), .B(data_point[29]), .Y(n25210) );
  INVXL U13577 ( .A(n22464), .Y(n22465) );
  NAND2XL U13578 ( .A(n23383), .B(n22463), .Y(n22466) );
  INVXL U13579 ( .A(n23038), .Y(n23044) );
  AOI211XL U13580 ( .A0(n23955), .A1(n23172), .B0(n23962), .C0(n23171), .Y(
        n25659) );
  INVXL U13581 ( .A(n23272), .Y(n23258) );
  INVXL U13582 ( .A(n23277), .Y(n23251) );
  AOI22XL U13583 ( .A0(n3017), .A1(n23177), .B0(n3040), .B1(n23176), .Y(n23191) );
  INVXL U13584 ( .A(n23175), .Y(n23192) );
  XOR2XL U13585 ( .A(n17182), .B(n17405), .Y(n17188) );
  ADDHXL U13586 ( .A(n25132), .B(n25131), .CO(n25133), .S(n25108) );
  INVXL U13587 ( .A(n23640), .Y(n23642) );
  AOI31XL U13588 ( .A0(n23788), .A1(n25699), .A2(n23787), .B0(n3115), .Y(
        n23791) );
  NAND2X1 U13589 ( .A(n5562), .B(n5401), .Y(n24425) );
  AOI21XL U13590 ( .A0(n23868), .A1(n23783), .B0(n23863), .Y(n5401) );
  NAND2X1 U13591 ( .A(n23864), .B(n23782), .Y(n5562) );
  NOR2X1 U13592 ( .A(n23780), .B(n23779), .Y(n24352) );
  INVXL U13593 ( .A(n23776), .Y(n23774) );
  INVXL U13594 ( .A(n23673), .Y(n23667) );
  NOR2X1 U13595 ( .A(n23666), .B(n23665), .Y(n25851) );
  XNOR2XL U13596 ( .A(n23663), .B(n23662), .Y(n23664) );
  NAND3X1 U13597 ( .A(n5568), .B(n5571), .C(n5570), .Y(n23839) );
  NAND2X1 U13598 ( .A(n23868), .B(n23686), .Y(n5570) );
  AOI22XL U13599 ( .A0(n25025), .A1(y12[17]), .B0(n3050), .B1(y11[17]), .Y(
        n24844) );
  AOI22XL U13600 ( .A0(n22486), .A1(sigma11[2]), .B0(n25754), .B1(sigma12[2]), 
        .Y(n20319) );
  NAND2X1 U13601 ( .A(n21048), .B(n5336), .Y(n5850) );
  AOI22XL U13602 ( .A0(n24739), .A1(y12[13]), .B0(n3050), .B1(y11[13]), .Y(
        n24704) );
  AOI22XL U13603 ( .A0(n24739), .A1(y12[9]), .B0(n25656), .B1(y11[9]), .Y(
        n24623) );
  AOI22XL U13604 ( .A0(n25025), .A1(y10[19]), .B0(n8104), .B1(y12[19]), .Y(
        n23834) );
  AOI22XL U13605 ( .A0(n24739), .A1(y12[10]), .B0(n3050), .B1(y11[10]), .Y(
        n24638) );
  AOI21XL U13606 ( .A0(n24824), .A1(n3060), .B0(n24823), .Y(n2425) );
  AOI22XL U13607 ( .A0(n25025), .A1(y12[16]), .B0(n25656), .B1(y11[16]), .Y(
        n24822) );
  AOI22XL U13608 ( .A0(n22486), .A1(sigma11[23]), .B0(sigma12[23]), .B1(n25754), .Y(n25811) );
  AOI22XL U13609 ( .A0(n22486), .A1(sigma11[26]), .B0(sigma12[26]), .B1(n25754), .Y(n25186) );
  AOI22XL U13610 ( .A0(n22486), .A1(sigma11[28]), .B0(sigma12[28]), .B1(n25754), .Y(n25164) );
  AOI22XL U13611 ( .A0(n25815), .A1(y10[6]), .B0(n25656), .B1(y12[6]), .Y(
        n24567) );
  AOI22XL U13612 ( .A0(n22486), .A1(sigma11[30]), .B0(sigma12[30]), .B1(n25754), .Y(n25794) );
  AOI22XL U13613 ( .A0(n25025), .A1(y10[18]), .B0(n8104), .B1(y12[18]), .Y(
        n23617) );
  AOI22XL U13614 ( .A0(n25815), .A1(y10[8]), .B0(n25656), .B1(y12[8]), .Y(
        n23584) );
  AOI22XL U13615 ( .A0(n25815), .A1(y12[4]), .B0(n3050), .B1(y11[4]), .Y(
        n24519) );
  AOI22XL U13616 ( .A0(n25815), .A1(y12[5]), .B0(n25656), .B1(y11[5]), .Y(
        n24542) );
  AOI21XL U13617 ( .A0(n4976), .A1(n21167), .B0(n21042), .Y(n2275) );
  AOI22XL U13618 ( .A0(n22486), .A1(sigma11[11]), .B0(n25754), .B1(sigma12[11]), .Y(n21041) );
  AOI22XL U13619 ( .A0(n25025), .A1(y10[20]), .B0(n3050), .B1(y12[20]), .Y(
        n23840) );
  AOI22XL U13620 ( .A0(n25815), .A1(y12[2]), .B0(n3050), .B1(y11[2]), .Y(
        n24485) );
  AOI22XL U13621 ( .A0(n25025), .A1(y12[1]), .B0(n3050), .B1(y11[1]), .Y(
        n24470) );
  OAI22XL U13622 ( .A0(n25255), .A1(n26138), .B0(n3050), .B1(n26414), .Y(
        n25192) );
  AOI22XL U13623 ( .A0(n25815), .A1(y12[26]), .B0(n3120), .B1(y11[26]), .Y(
        n25261) );
  OAI22XL U13624 ( .A0(n25754), .A1(n26137), .B0(n3059), .B1(n26416), .Y(
        n25200) );
  MXI2XL U13625 ( .A(mul5_out[29]), .B(n25209), .S0(n5770), .Y(n2354) );
  OAI21XL U13626 ( .A0(n24407), .A1(n3057), .B0(n24406), .Y(n24408) );
  AOI22XL U13627 ( .A0(n25025), .A1(y10[27]), .B0(n3050), .B1(y12[27]), .Y(
        n24406) );
  OAI21XL U13628 ( .A0(n25558), .A1(n25584), .B0(n25557), .Y(n2033) );
  AOI22XL U13629 ( .A0(n3051), .A1(n26127), .B0(n3061), .B1(n26478), .Y(n25557) );
  OAI21XL U13630 ( .A0(n25545), .A1(n3226), .B0(n25544), .Y(n2037) );
  AOI22XL U13631 ( .A0(n4575), .A1(n26126), .B0(n3061), .B1(n26477), .Y(n25544) );
  OAI21XL U13632 ( .A0(n25566), .A1(n4571), .B0(n25565), .Y(n2029) );
  AOI22XL U13633 ( .A0(n4575), .A1(n26128), .B0(n23088), .B1(n26479), .Y(
        n25565) );
  AOI22XL U13634 ( .A0(n3023), .A1(n26129), .B0(n23088), .B1(n26480), .Y(
        n25576) );
  AOI22XL U13635 ( .A0(n4575), .A1(n26111), .B0(n3061), .B1(n26459), .Y(n24371) );
  AOI22XL U13636 ( .A0(n3052), .A1(n26109), .B0(n3061), .B1(n26457), .Y(n24076) );
  AOI22XL U13637 ( .A0(n3052), .A1(n26110), .B0(n3061), .B1(n26458), .Y(n24320) );
  AOI22XL U13638 ( .A0(n4575), .A1(n26114), .B0(n3061), .B1(n26461), .Y(n25226) );
  AOI22XL U13639 ( .A0(n3052), .A1(n26112), .B0(n3061), .B1(n26486), .Y(n24457) );
  AOI22XL U13640 ( .A0(n3052), .A1(n26113), .B0(n3061), .B1(n26460), .Y(n25110) );
  AOI22XL U13641 ( .A0(n25410), .A1(n26134), .B0(n3061), .B1(n26485), .Y(
        n25800) );
  OAI21XL U13642 ( .A0(n23766), .A1(n3057), .B0(n23765), .Y(n23767) );
  AOI22XL U13643 ( .A0(n25815), .A1(y10[3]), .B0(n3050), .B1(y12[3]), .Y(
        n24511) );
  AOI22XL U13644 ( .A0(n25815), .A1(y10[7]), .B0(n25656), .B1(y12[7]), .Y(
        n23698) );
  AOI22XL U13645 ( .A0(n24739), .A1(y10[21]), .B0(n3050), .B1(y12[21]), .Y(
        n25029) );
  AOI22XL U13646 ( .A0(n22486), .A1(sigma11[1]), .B0(n25754), .B1(sigma12[1]), 
        .Y(n25295) );
  AOI22XL U13647 ( .A0(n22486), .A1(sigma11[14]), .B0(n25754), .B1(sigma12[14]), .Y(n24203) );
  AOI22XL U13648 ( .A0(n22486), .A1(sigma11[12]), .B0(n25754), .B1(sigma12[12]), .Y(n24185) );
  AOI22XL U13649 ( .A0(n22486), .A1(sigma11[5]), .B0(n25754), .B1(sigma12[5]), 
        .Y(n24137) );
  AOI22XL U13650 ( .A0(n22486), .A1(sigma11[4]), .B0(n25754), .B1(sigma12[4]), 
        .Y(n21025) );
  AOI22XL U13651 ( .A0(n22486), .A1(sigma11[10]), .B0(n25754), .B1(sigma12[10]), .Y(n24171) );
  AOI22XL U13652 ( .A0(n22486), .A1(sigma11[6]), .B0(n25754), .B1(sigma12[6]), 
        .Y(n21027) );
  AOI22XL U13653 ( .A0(n22486), .A1(sigma11[8]), .B0(n25754), .B1(sigma12[8]), 
        .Y(n21033) );
  AOI22XL U13654 ( .A0(n22486), .A1(sigma11[15]), .B0(n25754), .B1(sigma12[15]), .Y(n24212) );
  AOI22XL U13655 ( .A0(n22486), .A1(sigma11[16]), .B0(n25754), .B1(sigma12[16]), .Y(n24221) );
  AOI22XL U13656 ( .A0(n25201), .A1(sigma11[20]), .B0(n25754), .B1(sigma12[20]), .Y(n17460) );
  OAI21XL U13657 ( .A0(n24226), .A1(n5032), .B0(n24225), .Y(n5925) );
  AOI22XL U13658 ( .A0(n22486), .A1(sigma12[17]), .B0(n25750), .B1(sigma11[17]), .Y(n24225) );
  AOI22XL U13659 ( .A0(n22486), .A1(sigma11[18]), .B0(n25754), .B1(sigma12[18]), .Y(n24238) );
  AOI22XL U13660 ( .A0(n25201), .A1(sigma11[21]), .B0(n25754), .B1(sigma12[21]), .Y(n20842) );
  AOI21XL U13661 ( .A0(n5967), .A1(n21167), .B0(n21047), .Y(n2283) );
  AOI22XL U13662 ( .A0(n22486), .A1(sigma11[19]), .B0(n25754), .B1(sigma12[19]), .Y(n21046) );
  AOI22XL U13663 ( .A0(n25763), .A1(n26547), .B0(n25754), .B1(n26451), .Y(
        n25764) );
  OAI21XL U13664 ( .A0(n24157), .A1(n4875), .B0(n24156), .Y(n24158) );
  AOI22XL U13665 ( .A0(n22486), .A1(sigma12[9]), .B0(n25750), .B1(sigma11[9]), 
        .Y(n24156) );
  AOI22XL U13666 ( .A0(n25255), .A1(sigma12[2]), .B0(n3050), .B1(sigma11[2]), 
        .Y(n21053) );
  MXI2X1 U13667 ( .A(n24122), .B(n20749), .S0(n3111), .Y(n20750) );
  OAI21XL U13668 ( .A0(mul5_out[26]), .A1(n5015), .B0(n25182), .Y(n2348) );
  AOI22XL U13669 ( .A0(n25763), .A1(n6220), .B0(n25754), .B1(n26456), .Y(
        n25182) );
  OAI21XL U13670 ( .A0(mul5_out[28]), .A1(n4875), .B0(n25163), .Y(n2352) );
  AOI22XL U13671 ( .A0(n25786), .A1(n26106), .B0(n25785), .B1(n26452), .Y(
        n25163) );
  AOI22XL U13672 ( .A0(n25410), .A1(n26125), .B0(n3061), .B1(n26474), .Y(
        n25507) );
  OAI21XL U13673 ( .A0(n25485), .A1(n4573), .B0(n25484), .Y(n2057) );
  AOI22XL U13674 ( .A0(n3052), .A1(n26136), .B0(n3061), .B1(n26472), .Y(n25484) );
  OAI21XL U13675 ( .A0(n25459), .A1(n3226), .B0(n25458), .Y(n2065) );
  AOI22XL U13676 ( .A0(n3052), .A1(n26122), .B0(n3061), .B1(n26470), .Y(n25458) );
  OAI21XL U13677 ( .A0(n25371), .A1(n3226), .B0(n25370), .Y(n2093) );
  AOI22XL U13678 ( .A0(n4575), .A1(n26116), .B0(n3061), .B1(n26463), .Y(n25370) );
  OAI2BB1XL U13679 ( .A0N(w1[352]), .A1N(n3052), .B0(n25645), .Y(n25646) );
  AOI22XL U13680 ( .A0(n3028), .A1(w1[256]), .B0(in_valid_w1), .B1(weight1[0]), 
        .Y(n25645) );
  OAI2BB1XL U13681 ( .A0N(w1[356]), .A1N(n25410), .B0(n25580), .Y(n25581) );
  AOI22XL U13682 ( .A0(n3064), .A1(w1[260]), .B0(in_valid_w1), .B1(weight1[4]), 
        .Y(n25580) );
  OAI2BB1XL U13683 ( .A0N(w1[374]), .A1N(n25410), .B0(n25365), .Y(n25366) );
  AOI22XL U13684 ( .A0(n3028), .A1(w1[278]), .B0(in_valid_w1), .B1(weight1[22]), .Y(n25365) );
  OAI2BB2XL U13685 ( .B0(n22903), .B1(n3225), .A0N(n22987), .A1N(n22904), .Y(
        n10807) );
  NAND2XL U13686 ( .A(n22932), .B(n22987), .Y(n4709) );
  OAI2BB2XL U13687 ( .B0(n22981), .B1(n3225), .A0N(n22987), .A1N(n22980), .Y(
        n22982) );
  XOR2XL U13688 ( .A(n22991), .B(n22990), .Y(n23000) );
  NAND2XL U13689 ( .A(n22988), .B(n22987), .Y(n4705) );
  NAND2BXL U13690 ( .AN(n3110), .B(n3211), .Y(n16397) );
  XNOR2XL U13691 ( .A(n25869), .B(n25878), .Y(n7066) );
  INVXL U13692 ( .A(n15281), .Y(n15089) );
  XNOR2X1 U13693 ( .A(M2_mult_x_15_a_1_), .B(n10311), .Y(n9962) );
  OAI22XL U13694 ( .A0(n12357), .A1(n12285), .B0(n12284), .B1(n12283), .Y(
        n12287) );
  NAND2BXL U13695 ( .AN(n3110), .B(n12282), .Y(n12283) );
  OAI22XL U13696 ( .A0(n12340), .A1(M3_mult_x_15_b_1_), .B0(n12280), .B1(
        n12338), .Y(n12275) );
  NOR2BXL U13697 ( .AN(n3110), .B(n12284), .Y(n12274) );
  NAND2BXL U13698 ( .AN(n3110), .B(n2980), .Y(n12272) );
  XNOR2XL U13699 ( .A(n12233), .B(n11499), .Y(n12350) );
  XNOR2X1 U13700 ( .A(n2980), .B(n3021), .Y(n12064) );
  XNOR2XL U13701 ( .A(n14028), .B(n13605), .Y(n13075) );
  INVXL U13702 ( .A(n8557), .Y(n8238) );
  INVXL U13703 ( .A(n8552), .Y(n8319) );
  INVXL U13704 ( .A(n8534), .Y(n8342) );
  INVXL U13705 ( .A(n8532), .Y(n8340) );
  INVXL U13706 ( .A(n19625), .Y(n19472) );
  INVXL U13707 ( .A(n19623), .Y(n19470) );
  INVXL U13708 ( .A(n19646), .Y(n19368) );
  INVXL U13709 ( .A(n15320), .Y(n14984) );
  INVXL U13710 ( .A(n21691), .Y(n21644) );
  INVXL U13711 ( .A(n15351), .Y(n15247) );
  INVXL U13712 ( .A(n15296), .Y(n15193) );
  INVXL U13713 ( .A(n15334), .Y(n15079) );
  INVXL U13714 ( .A(n21676), .Y(n21544) );
  INVXL U13715 ( .A(n21717), .Y(n21539) );
  NAND2XL U13716 ( .A(n21689), .B(n21537), .Y(n21538) );
  INVXL U13717 ( .A(n21731), .Y(n21537) );
  NAND2XL U13718 ( .A(n21643), .B(n21532), .Y(n21533) );
  INVXL U13719 ( .A(n21698), .Y(n21532) );
  XOR2XL U13720 ( .A(n22973), .B(n3055), .Y(n23020) );
  XOR2XL U13721 ( .A(n22979), .B(n3056), .Y(n23029) );
  AOI222XL U13722 ( .A0(n22988), .A1(n10749), .B0(n22980), .B1(n3116), .C0(
        n22976), .C1(n22987), .Y(n22977) );
  NOR2BX1 U13723 ( .AN(n6944), .B(n7634), .Y(n6396) );
  NAND2BXL U13724 ( .AN(n6944), .B(n25869), .Y(n6398) );
  XNOR2XL U13725 ( .A(n4806), .B(n23220), .Y(n6425) );
  XNOR2XL U13726 ( .A(n4806), .B(n25866), .Y(n6555) );
  XNOR2XL U13727 ( .A(n4806), .B(n21054), .Y(n6572) );
  XNOR2XL U13728 ( .A(M0_b_1_), .B(n25866), .Y(n6571) );
  OAI22XL U13729 ( .A0(n6573), .A1(n6845), .B0(n6572), .B1(n6843), .Y(n6574)
         );
  XNOR2XL U13730 ( .A(M0_b_1_), .B(n3209), .Y(n6554) );
  XNOR2XL U13731 ( .A(n25866), .B(n7165), .Y(n6603) );
  XNOR2XL U13732 ( .A(n25866), .B(n7164), .Y(n6601) );
  XNOR2XL U13733 ( .A(M0_b_1_), .B(n25867), .Y(n6614) );
  XNOR2XL U13734 ( .A(n4806), .B(n25867), .Y(n6515) );
  NAND2BXL U13735 ( .AN(n6944), .B(n23220), .Y(n6460) );
  XNOR2XL U13736 ( .A(M0_b_1_), .B(n23221), .Y(n6330) );
  OAI21X2 U13737 ( .A0(n7382), .A1(n26006), .B0(n6236), .Y(M0_a_3_) );
  OAI21XL U13738 ( .A0(n7382), .A1(n26009), .B0(n6230), .Y(M0_a_0_) );
  AOI21XL U13739 ( .A0(n6733), .A1(y10[0]), .B0(n24266), .Y(n6230) );
  INVXL U13740 ( .A(n10850), .Y(n10851) );
  OAI22XL U13741 ( .A0(n16638), .A1(n2978), .B0(M3_mult_x_15_b_1_), .B1(n16475), .Y(n16622) );
  XNOR2XL U13742 ( .A(M5_mult_x_15_n1), .B(n11499), .Y(n16636) );
  XNOR2XL U13743 ( .A(n3047), .B(n12271), .Y(n16639) );
  XNOR2XL U13744 ( .A(n3047), .B(M3_mult_x_15_b_1_), .Y(n16640) );
  NAND2BXL U13745 ( .AN(n16639), .B(n5847), .Y(n5839) );
  CMPR32X1 U13746 ( .A(n16608), .B(n16607), .C(n16606), .CO(n16600), .S(n16610) );
  OAI22XL U13747 ( .A0(n16701), .A1(n16615), .B0(n16699), .B1(n16594), .Y(
        n16606) );
  CMPR32X1 U13748 ( .A(n16597), .B(n16596), .C(n16595), .CO(n16589), .S(n16599) );
  OAI22XL U13749 ( .A0(n16701), .A1(n16594), .B0(n16699), .B1(n16584), .Y(
        n16595) );
  OAI22XL U13750 ( .A0(n3102), .A1(n16583), .B0(n16332), .B1(n16582), .Y(
        n16596) );
  NAND2BXL U13751 ( .AN(n3110), .B(n16289), .Y(n16571) );
  XNOR2XL U13752 ( .A(n3047), .B(M3_mult_x_15_b_6_), .Y(n16573) );
  NOR2BXL U13753 ( .AN(n3110), .B(n16688), .Y(n16580) );
  NAND2BXL U13754 ( .AN(n3110), .B(n15968), .Y(n16574) );
  NAND2BXL U13755 ( .AN(n16540), .B(n3044), .Y(n5844) );
  XOR2X1 U13756 ( .A(n15968), .B(M3_mult_x_15_b_3_), .Y(n5734) );
  NAND2BXL U13757 ( .AN(n3110), .B(n3203), .Y(n16517) );
  XNOR2XL U13758 ( .A(n15968), .B(n11499), .Y(n16516) );
  XOR2XL U13759 ( .A(n16614), .B(n16965), .Y(n16533) );
  XNOR2XL U13760 ( .A(n16614), .B(M3_mult_x_15_b_9_), .Y(n16498) );
  NAND2BXL U13761 ( .AN(n16408), .B(n3044), .Y(n5845) );
  XOR2XL U13762 ( .A(n16289), .B(n16965), .Y(n16474) );
  XNOR2XL U13763 ( .A(n16614), .B(M3_mult_x_15_b_13_), .Y(n16361) );
  XNOR2XL U13764 ( .A(n3203), .B(M3_mult_x_15_b_6_), .Y(n16346) );
  XNOR2XL U13765 ( .A(n3047), .B(n11495), .Y(n16381) );
  NAND2XL U13766 ( .A(n10772), .B(n10771), .Y(n10811) );
  NOR2XL U13767 ( .A(n26496), .B(n10775), .Y(n10854) );
  NOR2XL U13768 ( .A(n10769), .B(n10775), .Y(n10788) );
  NAND2XL U13769 ( .A(n26496), .B(n10775), .Y(n10855) );
  OAI2BB1XL U13770 ( .A0N(n7060), .A1N(n7059), .B0(n7058), .Y(n7067) );
  OAI21XL U13771 ( .A0(n7053), .A1(n7695), .B0(n5120), .Y(n7069) );
  NAND2XL U13772 ( .A(n7057), .B(M0_b_1_), .Y(n7058) );
  NOR2XL U13773 ( .A(n6861), .B(n6843), .Y(n6943) );
  XNOR2XL U13774 ( .A(n25869), .B(n25880), .Y(n6924) );
  NAND2X1 U13775 ( .A(n5114), .B(n5113), .Y(n7030) );
  XNOR2X1 U13776 ( .A(n7057), .B(n7056), .Y(n6992) );
  NAND2BXL U13777 ( .AN(n7184), .B(n5122), .Y(n5115) );
  CLKINVX3 U13778 ( .A(M2_a_7_), .Y(n9201) );
  OAI22XL U13779 ( .A0(n9983), .A1(n9907), .B0(n9906), .B1(n9905), .Y(n9909)
         );
  OAI22XL U13780 ( .A0(n9963), .A1(n9960), .B0(n3182), .B1(n3180), .Y(n9895)
         );
  NAND2BXL U13781 ( .AN(n9960), .B(M2_mult_x_15_a_1_), .Y(n9893) );
  NOR2BXL U13782 ( .AN(n9960), .B(n9981), .Y(n9896) );
  XNOR2X1 U13783 ( .A(n9904), .B(n9901), .Y(n9885) );
  OAI22XL U13784 ( .A0(n9979), .A1(n9878), .B0(n9977), .B1(n9876), .Y(n9889)
         );
  NAND2BXL U13785 ( .AN(n9960), .B(n9886), .Y(n9876) );
  ADDFX2 U13786 ( .A(n9881), .B(n9880), .CI(n9879), .CO(n9871), .S(n9882) );
  OAI22XL U13787 ( .A0(n9979), .A1(n9887), .B0(n9977), .B1(n9865), .Y(n9879)
         );
  OAI22XL U13788 ( .A0(n9963), .A1(n9875), .B0(n9864), .B1(n3180), .Y(n9880)
         );
  OAI22XL U13789 ( .A0(n9979), .A1(n9865), .B0(n9977), .B1(n9854), .Y(n9866)
         );
  NOR2BXL U13790 ( .AN(n9960), .B(n10159), .Y(n9849) );
  XNOR2XL U13791 ( .A(n9904), .B(n10312), .Y(n9980) );
  NOR2X1 U13792 ( .A(n9087), .B(n25902), .Y(n5348) );
  NAND2X1 U13793 ( .A(n9164), .B(target_temp[5]), .Y(n11531) );
  AOI22XL U13794 ( .A0(n11536), .A1(data[3]), .B0(in_valid_d), .B1(w1[259]), 
        .Y(n9101) );
  NOR2X1 U13795 ( .A(n25243), .B(n23999), .Y(n5090) );
  XNOR2XL U13796 ( .A(M2_a_17_), .B(n10311), .Y(n9208) );
  NOR2BXL U13797 ( .AN(n3110), .B(n12595), .Y(n12349) );
  CMPR32X1 U13798 ( .A(n12346), .B(n12345), .C(n12344), .CO(n12367), .S(n12375) );
  CMPR32X1 U13799 ( .A(n12231), .B(n12230), .C(n12229), .CO(n12364), .S(n12242) );
  NOR2BXL U13800 ( .AN(n3110), .B(n12342), .Y(n12231) );
  NAND2BXL U13801 ( .AN(n3110), .B(n12233), .Y(n12221) );
  OAI22XL U13802 ( .A0(n12152), .A1(n12246), .B0(n3185), .B1(n12236), .Y(
        n12247) );
  ADDFX2 U13803 ( .A(n12263), .B(n4800), .CI(n12261), .CO(n12316), .S(n12315)
         );
  OAI22XL U13804 ( .A0(n12357), .A1(n12264), .B0(n12284), .B1(n12254), .Y(
        n12263) );
  ADDHXL U13805 ( .A(n12297), .B(n12296), .CO(n12298), .S(n12288) );
  OAI22XL U13806 ( .A0(n12357), .A1(n12281), .B0(n12284), .B1(n12295), .Y(
        n12296) );
  OAI22XL U13807 ( .A0(n12340), .A1(n12280), .B0(n12292), .B1(n12338), .Y(
        n12297) );
  OAI22XL U13808 ( .A0(n12357), .A1(n12295), .B0(n12284), .B1(n12294), .Y(
        n12306) );
  OAI22XL U13809 ( .A0(n12293), .A1(n12292), .B0(n12291), .B1(n12338), .Y(
        n12307) );
  OAI22XL U13810 ( .A0(n12357), .A1(n12294), .B0(n12284), .B1(n12264), .Y(
        n12305) );
  NAND2BXL U13811 ( .AN(n3110), .B(n12594), .Y(n12187) );
  XOR2XL U13812 ( .A(n3108), .B(n12594), .Y(n6104) );
  XNOR2X1 U13813 ( .A(n12282), .B(n3190), .Y(n12150) );
  NOR2X1 U13814 ( .A(n5784), .B(n5783), .Y(n5782) );
  NOR2X1 U13815 ( .A(n5516), .B(n12597), .Y(n5784) );
  NOR2XL U13816 ( .A(n12001), .B(n12595), .Y(n5783) );
  XNOR2XL U13817 ( .A(n13769), .B(M1_b_3_), .Y(n13116) );
  XNOR2XL U13818 ( .A(n13919), .B(n13204), .Y(n13092) );
  OAI22XL U13819 ( .A0(n13116), .A1(n13721), .B0(n13108), .B1(n13790), .Y(
        n13110) );
  XNOR2XL U13820 ( .A(n13049), .B(M1_b_3_), .Y(n13108) );
  NOR2BXL U13821 ( .AN(n13049), .B(n13721), .Y(n13101) );
  NAND2BXL U13822 ( .AN(n13049), .B(n13605), .Y(n13098) );
  NOR2BXL U13823 ( .AN(n13049), .B(n14029), .Y(n13061) );
  OAI22XL U13824 ( .A0(n13065), .A1(n13721), .B0(n13074), .B1(n13790), .Y(
        n13076) );
  OAI22XL U13825 ( .A0(n14044), .A1(n6210), .B0(n13052), .B1(n13974), .Y(
        n13159) );
  NAND2BXL U13826 ( .AN(n13049), .B(n14030), .Y(n13052) );
  XOR2XL U13827 ( .A(n25865), .B(n5512), .Y(n13359) );
  INVXL U13828 ( .A(n4807), .Y(n13047) );
  XNOR2XL U13829 ( .A(n14195), .B(n25863), .Y(n14025) );
  XNOR2XL U13830 ( .A(n14236), .B(n25863), .Y(n14059) );
  CMPR32X1 U13831 ( .A(n14092), .B(n14091), .C(n14090), .CO(n14123), .S(n14101) );
  INVXL U13832 ( .A(n14118), .Y(n14092) );
  XNOR2X1 U13833 ( .A(n18006), .B(n3198), .Y(n17963) );
  OAI22XL U13834 ( .A0(n18239), .A1(n18130), .B0(n18238), .B1(n18120), .Y(
        n18131) );
  NOR2BXL U13835 ( .AN(n2978), .B(n18429), .Y(n18233) );
  OAI22XL U13836 ( .A0(n18111), .A1(n6096), .B0(n18227), .B1(n18504), .Y(
        n18231) );
  NAND2BXL U13837 ( .AN(n2978), .B(n18118), .Y(n18105) );
  OAI22XL U13838 ( .A0(n18107), .A1(n6036), .B0(n18113), .B1(n18235), .Y(
        n18114) );
  XNOR2X1 U13839 ( .A(n18150), .B(n3190), .Y(n17992) );
  XNOR2XL U13840 ( .A(n18503), .B(n11499), .Y(n18066) );
  XNOR2XL U13841 ( .A(n14028), .B(M1_b_19_), .Y(n13690) );
  OAI22XL U13842 ( .A0(n8467), .A1(n3087), .B0(n3157), .B1(n8484), .Y(n8468)
         );
  AOI21XL U13843 ( .A0(n3154), .A1(n8602), .B0(n8396), .Y(n8397) );
  AOI21XL U13844 ( .A0(n19807), .A1(n19687), .B0(n19527), .Y(n19528) );
  AOI2BB2XL U13845 ( .B0(n19501), .B1(n19542), .A0N(n19542), .A1N(n19711), .Y(
        n19601) );
  AOI2BB2XL U13846 ( .B0(n19709), .B1(n3036), .A0N(n3036), .A1N(n19708), .Y(
        n19710) );
  NAND2XL U13847 ( .A(n3041), .B(n19432), .Y(n19433) );
  NAND2XL U13848 ( .A(n3041), .B(n19442), .Y(n19443) );
  NAND2XL U13849 ( .A(n3041), .B(n19428), .Y(n19429) );
  INVXL U13850 ( .A(n19556), .Y(n19599) );
  INVXL U13851 ( .A(n19560), .Y(n19721) );
  INVXL U13852 ( .A(n19567), .Y(n19753) );
  INVXL U13853 ( .A(n19562), .Y(n19737) );
  INVXL U13854 ( .A(n19486), .Y(n19533) );
  INVXL U13855 ( .A(n19383), .Y(n19456) );
  NAND2XL U13856 ( .A(n15190), .B(n15063), .Y(n15064) );
  NAND2XL U13857 ( .A(n15190), .B(n15053), .Y(n15054) );
  NAND2XL U13858 ( .A(n15190), .B(n15050), .Y(n15051) );
  AOI2BB2XL U13859 ( .B0(n15190), .B1(n15048), .A0N(n15558), .A1N(n15548), .Y(
        n15281) );
  INVXL U13860 ( .A(n21743), .Y(n21645) );
  INVXL U13861 ( .A(n15227), .Y(n15260) );
  NAND2XL U13862 ( .A(n15215), .B(n15313), .Y(n15216) );
  AOI22XL U13863 ( .A0(n15232), .A1(n6194), .B0(n15214), .B1(n3016), .Y(n15215) );
  INVXL U13864 ( .A(n15213), .Y(n15214) );
  INVXL U13865 ( .A(n15544), .Y(n15218) );
  INVXL U13866 ( .A(n15174), .Y(n15207) );
  AOI2BB2XL U13867 ( .B0(n15265), .B1(n3156), .A0N(n3156), .A1N(n15179), .Y(
        n15180) );
  AOI22XL U13868 ( .A0(n15289), .A1(n15230), .B0(n3038), .B1(n15229), .Y(
        n15264) );
  INVXL U13869 ( .A(n15302), .Y(n15077) );
  INVXL U13870 ( .A(n15323), .Y(n15084) );
  INVXL U13871 ( .A(n15338), .Y(n15082) );
  INVXL U13872 ( .A(n15023), .Y(n15019) );
  NAND2XL U13873 ( .A(n15026), .B(n15033), .Y(n15028) );
  INVXL U13874 ( .A(n15033), .Y(n15034) );
  INVXL U13875 ( .A(n14995), .Y(n15076) );
  NAND2XL U13876 ( .A(n21847), .B(n3171), .Y(n21784) );
  NAND2XL U13877 ( .A(n21799), .B(n3037), .Y(n21800) );
  INVXL U13878 ( .A(n21796), .Y(n21797) );
  INVXL U13879 ( .A(n21984), .Y(n21804) );
  NAND2XL U13880 ( .A(n21580), .B(n21568), .Y(n21569) );
  INVXL U13881 ( .A(n21567), .Y(n21568) );
  AOI22XL U13882 ( .A0(n3095), .A1(n21563), .B0(n21562), .B1(n21580), .Y(
        n21767) );
  INVXL U13883 ( .A(n21561), .Y(n21562) );
  AOI22XL U13884 ( .A0(n3095), .A1(n21746), .B0(n21745), .B1(n21580), .Y(
        n21778) );
  INVXL U13885 ( .A(n21583), .Y(n21584) );
  NAND2XL U13886 ( .A(n21580), .B(n21524), .Y(n21525) );
  INVXL U13887 ( .A(n21566), .Y(n21524) );
  NAND2XL U13888 ( .A(n21580), .B(n21464), .Y(n21465) );
  INVXL U13889 ( .A(n21570), .Y(n21464) );
  AOI21XL U13890 ( .A0(n8517), .A1(n8601), .B0(n8610), .Y(n8374) );
  NAND2XL U13891 ( .A(n8512), .B(n3154), .Y(n8373) );
  NAND2XL U13892 ( .A(n8415), .B(n8593), .Y(n8416) );
  NAND2XL U13893 ( .A(n8413), .B(n3086), .Y(n8414) );
  AOI22XL U13894 ( .A0(n8499), .A1(n3087), .B0(n8412), .B1(n3157), .Y(n8413)
         );
  INVXL U13895 ( .A(n23003), .Y(n22970) );
  AOI222XL U13896 ( .A0(n23152), .A1(n11058), .B0(n23093), .B1(n23151), .C0(
        n23150), .C1(n10789), .Y(n23141) );
  INVXL U13897 ( .A(n23023), .Y(n22886) );
  XOR2X1 U13898 ( .A(n7139), .B(n7141), .Y(n5105) );
  XOR2XL U13899 ( .A(n22704), .B(n3058), .Y(n23037) );
  INVXL U13900 ( .A(n22702), .Y(n22703) );
  AOI222XL U13901 ( .A0(n22988), .A1(n10775), .B0(n22980), .B1(n10769), .C0(
        n22976), .C1(n23002), .Y(n22743) );
  AOI222XL U13902 ( .A0(n23003), .A1(n23151), .B0(n22969), .B1(n10789), .C0(
        n23001), .C1(n3220), .Y(n21088) );
  AOI222XL U13903 ( .A0(n22988), .A1(n26496), .B0(n22980), .B1(n10775), .C0(
        n22976), .C1(n10769), .Y(n22921) );
  XOR2XL U13904 ( .A(n22798), .B(n3221), .Y(M6_mult_x_15_n1204) );
  NOR2XL U13905 ( .A(n26493), .B(n11059), .Y(n22763) );
  INVXL U13906 ( .A(n22759), .Y(n22760) );
  XOR2XL U13907 ( .A(n22724), .B(n3058), .Y(n23034) );
  AOI222XL U13908 ( .A0(n22928), .A1(n23002), .B0(n22700), .B1(n10749), .C0(
        n22927), .C1(n3116), .Y(n22723) );
  AOI222XL U13909 ( .A0(n23003), .A1(n11058), .B0(n22969), .B1(n23151), .C0(
        n23001), .C1(n10789), .Y(n22937) );
  AOI222XL U13910 ( .A0(n22988), .A1(n3220), .B0(n22980), .B1(n22867), .C0(
        n22976), .C1(n10775), .Y(n22847) );
  XOR2XL U13911 ( .A(n23027), .B(n3054), .Y(M6_mult_x_15_n1149) );
  AOI222XL U13912 ( .A0(n23023), .A1(n3217), .B0(n22887), .B1(n23022), .C0(
        n23021), .C1(n11059), .Y(n23024) );
  NOR2XL U13913 ( .A(n11058), .B(n23151), .Y(n22644) );
  NAND2XL U13914 ( .A(n11058), .B(n23151), .Y(n22645) );
  AOI21XL U13915 ( .A0(n22587), .A1(n22586), .B0(n22585), .Y(n22588) );
  NAND2XL U13916 ( .A(n22583), .B(n22586), .Y(n22589) );
  INVXL U13917 ( .A(n22584), .Y(n22587) );
  INVXL U13918 ( .A(n22590), .Y(n22630) );
  INVXL U13919 ( .A(n22629), .Y(n22591) );
  NAND2XL U13920 ( .A(n26493), .B(n3217), .Y(n22772) );
  XNOR2XL U13921 ( .A(n10825), .B(n10824), .Y(n23006) );
  NAND2XL U13922 ( .A(n10823), .B(n10822), .Y(n10825) );
  INVXL U13923 ( .A(n11139), .Y(n10823) );
  XOR2XL U13924 ( .A(n22712), .B(n3119), .Y(n22719) );
  INVXL U13925 ( .A(n22710), .Y(n22711) );
  NAND2XL U13926 ( .A(n3116), .B(n10749), .Y(n10772) );
  NAND2XL U13927 ( .A(n3116), .B(n22987), .Y(n10771) );
  NAND2XL U13928 ( .A(n10769), .B(n10775), .Y(n10850) );
  INVXL U13929 ( .A(n11056), .Y(n10853) );
  INVXL U13930 ( .A(n10788), .Y(n10852) );
  INVXL U13931 ( .A(n22602), .Y(n22603) );
  INVXL U13932 ( .A(n22601), .Y(n22604) );
  INVXL U13933 ( .A(n22605), .Y(n22761) );
  XNOR2XL U13934 ( .A(n21063), .B(n21062), .Y(n21064) );
  XNOR2XL U13935 ( .A(n3055), .B(n21062), .Y(n22563) );
  XOR2XL U13936 ( .A(n3056), .B(n21063), .Y(n22562) );
  NAND2XL U13937 ( .A(n11063), .B(n11073), .Y(n22567) );
  INVXL U13938 ( .A(n22575), .Y(n22774) );
  INVXL U13939 ( .A(n22772), .Y(n22773) );
  NAND2XL U13940 ( .A(n11062), .B(n3217), .Y(n22777) );
  XNOR2XL U13941 ( .A(n25869), .B(n6944), .Y(n6409) );
  OAI22XL U13942 ( .A0(M0_b_1_), .A1(n6845), .B0(n6573), .B1(n6843), .Y(n6568)
         );
  OAI22XL U13943 ( .A0(n6616), .A1(n7093), .B0(n6615), .B1(n7094), .Y(n6625)
         );
  CMPR32X1 U13944 ( .A(n6645), .B(n6644), .C(n6643), .CO(n6518), .S(n6654) );
  OAI22XL U13945 ( .A0(n6501), .A1(n6843), .B0(n6845), .B1(n6516), .Y(n6644)
         );
  OAI2BB1XL U13946 ( .A0N(n5631), .A1N(n6498), .B0(n5630), .Y(n6506) );
  NAND2XL U13947 ( .A(n5634), .B(n6499), .Y(n5630) );
  NAND2BXL U13948 ( .AN(n5634), .B(n5632), .Y(n5631) );
  XNOR2XL U13949 ( .A(n3209), .B(n25880), .Y(n6449) );
  CLKINVX2 U13950 ( .A(n6366), .Y(n6602) );
  OAI22XL U13951 ( .A0(n7633), .A1(n7615), .B0(n7634), .B1(n6320), .Y(n6375)
         );
  NAND2BXL U13952 ( .AN(n6944), .B(n23221), .Y(n6320) );
  CMPR32X1 U13953 ( .A(n6318), .B(n6317), .C(n6316), .CO(n6334), .S(n6372) );
  OAI22XL U13954 ( .A0(n6327), .A1(n4592), .B0(n3046), .B1(n6314), .Y(n6318)
         );
  OAI21XL U13955 ( .A0(n7828), .A1(n6944), .B0(n7829), .Y(n6860) );
  XNOR2X1 U13956 ( .A(n3209), .B(n7646), .Y(n6780) );
  XNOR2X1 U13957 ( .A(n21054), .B(n25874), .Y(n6290) );
  INVX1 U13958 ( .A(M0_a_6_), .Y(n5628) );
  INVXL U13959 ( .A(n21085), .Y(n22643) );
  NAND2XL U13960 ( .A(n10789), .B(n23151), .Y(n22641) );
  INVXL U13961 ( .A(n22932), .Y(n22903) );
  NOR2XL U13962 ( .A(n10789), .B(n3220), .Y(n11046) );
  AOI21XL U13963 ( .A0(n10853), .A1(n11048), .B0(n11052), .Y(n10872) );
  NOR2XL U13964 ( .A(n26496), .B(n3220), .Y(n11047) );
  OAI22XL U13965 ( .A0(n16942), .A1(n16467), .B0(n16688), .B1(n16401), .Y(
        n16472) );
  OAI22XL U13966 ( .A0(n16701), .A1(n16700), .B0(n16699), .B1(n16698), .Y(
        n16709) );
  CMPR32X1 U13967 ( .A(n16692), .B(n16691), .C(n16690), .CO(n16714), .S(n16722) );
  OAI22XL U13968 ( .A0(n16942), .A1(n16568), .B0(n16688), .B1(n16689), .Y(
        n16691) );
  CMPR32X1 U13969 ( .A(n16501), .B(n16500), .C(n16499), .CO(n16551), .S(n16507) );
  NAND2BXL U13970 ( .AN(n3110), .B(n3199), .Y(n16477) );
  OAI22XL U13971 ( .A0(n16701), .A1(n16473), .B0(n16699), .B1(n16459), .Y(
        n16492) );
  XNOR2XL U13972 ( .A(n16289), .B(n3190), .Y(n16351) );
  NAND2BXL U13973 ( .AN(n3110), .B(n17039), .Y(n16334) );
  XNOR2X1 U13974 ( .A(n3199), .B(n3190), .Y(n16002) );
  NAND2BXL U13975 ( .AN(n3110), .B(n17073), .Y(n16109) );
  OAI22XL U13976 ( .A0(n17060), .A1(n5704), .B0(n16377), .B1(n17061), .Y(
        n16338) );
  NAND2XL U13977 ( .A(learning_rate[3]), .B(in_valid_t), .Y(n4754) );
  AOI2BB1XL U13978 ( .A0N(n11146), .A1N(n11145), .B0(n11144), .Y(n11148) );
  AOI2BB1XL U13979 ( .A0N(n11143), .A1N(n11142), .B0(n11141), .Y(n11145) );
  AOI21XL U13980 ( .A0(n10774), .A1(n10811), .B0(n10773), .Y(n11056) );
  NOR2XL U13981 ( .A(n10812), .B(n11139), .Y(n10774) );
  NAND2XL U13982 ( .A(n10813), .B(n10822), .Y(n10773) );
  NOR2XL U13983 ( .A(n10788), .B(n10854), .Y(n11048) );
  NOR2XL U13984 ( .A(n11047), .B(n11046), .Y(n11053) );
  NAND2XL U13985 ( .A(n10855), .B(n10850), .Y(n11052) );
  NAND2XL U13986 ( .A(n26496), .B(n3220), .Y(n11049) );
  NAND2XL U13987 ( .A(n10789), .B(n3220), .Y(n11050) );
  NOR2XL U13988 ( .A(n22642), .B(n22644), .Y(n22601) );
  NOR2XL U13989 ( .A(n26493), .B(n3217), .Y(n22575) );
  NOR2XL U13990 ( .A(n11062), .B(n3217), .Y(n22776) );
  NOR2XL U13991 ( .A(n11062), .B(n23109), .Y(n22590) );
  NOR2XL U13992 ( .A(n11063), .B(n23109), .Y(n22592) );
  NAND2XL U13993 ( .A(n22777), .B(n22772), .Y(n22585) );
  NAND2XL U13994 ( .A(n11063), .B(n23109), .Y(n22593) );
  NAND2XL U13995 ( .A(n11062), .B(n23109), .Y(n22629) );
  NAND2XL U13996 ( .A(n22645), .B(n22641), .Y(n22602) );
  NAND2XL U13997 ( .A(n26493), .B(n11059), .Y(n22764) );
  NAND2XL U13998 ( .A(n11058), .B(n11059), .Y(n22759) );
  NOR2XL U13999 ( .A(n22605), .B(n22763), .Y(n11061) );
  NOR2XL U14000 ( .A(n22553), .B(n22555), .Y(n22496) );
  NAND2XL U14001 ( .A(n22556), .B(n22567), .Y(n22497) );
  NOR2XL U14002 ( .A(n22500), .B(n22530), .Y(n11076) );
  XNOR2X1 U14003 ( .A(n17038), .B(n3043), .Y(n16938) );
  INVXL U14004 ( .A(n8253), .Y(n8327) );
  NAND2XL U14005 ( .A(n8482), .B(n8303), .Y(n8304) );
  NAND2XL U14006 ( .A(n8482), .B(n8299), .Y(n8300) );
  INVXL U14007 ( .A(n8479), .Y(n8510) );
  NAND2XL U14008 ( .A(n3040), .B(n8256), .Y(n8257) );
  INVXL U14009 ( .A(n8422), .Y(n8444) );
  INVXL U14010 ( .A(n8354), .Y(n8379) );
  INVXL U14011 ( .A(n8427), .Y(n8475) );
  XNOR2X1 U14012 ( .A(n8227), .B(n8226), .Y(n8537) );
  OR2X2 U14013 ( .A(n6833), .B(n7094), .Y(n5129) );
  XNOR2XL U14014 ( .A(n4806), .B(n23219), .Y(n6847) );
  XNOR2XL U14015 ( .A(n25866), .B(n7800), .Y(n6834) );
  OAI22XL U14016 ( .A0(n7093), .A1(n6963), .B0(n7027), .B1(n3599), .Y(n7034)
         );
  OAI22X1 U14017 ( .A0(n7829), .A1(n4806), .B0(n7828), .B1(n7165), .Y(n7037)
         );
  CMPR32X1 U14018 ( .A(n7158), .B(n7157), .C(n7156), .CO(n7179), .S(n7155) );
  OAI21XL U14019 ( .A0(n7695), .A1(n7148), .B0(n5116), .Y(n7156) );
  OAI22XL U14020 ( .A0(n7633), .A1(n7197), .B0(n7232), .B1(n6300), .Y(n7235)
         );
  OAI22XL U14021 ( .A0(n7535), .A1(n7291), .B0(n7461), .B1(n7460), .Y(n7464)
         );
  CMPR32X1 U14022 ( .A(n7285), .B(n7284), .C(n7283), .CO(n7470), .S(n7281) );
  OAI22XL U14023 ( .A0(n7511), .A1(n7221), .B0(n7512), .B1(n7289), .Y(n7284)
         );
  OAI21X1 U14024 ( .A0(n7227), .A1(n7695), .B0(n5117), .Y(n7217) );
  XNOR2XL U14025 ( .A(n25885), .B(n10311), .Y(n9506) );
  XNOR2X1 U14026 ( .A(M2_a_17_), .B(n10386), .Y(n9505) );
  CMPR32X1 U14027 ( .A(n9339), .B(n9338), .C(n9337), .CO(n9476), .S(n9331) );
  OAI22XL U14028 ( .A0(n9590), .A1(n9219), .B0(n9877), .B1(n9886), .Y(n9338)
         );
  CMPR32X1 U14029 ( .A(n10156), .B(n10155), .C(n10154), .CO(n10304), .S(n10152) );
  NAND2X1 U14030 ( .A(n6059), .B(n9841), .Y(n10297) );
  INVXL U14031 ( .A(n10342), .Y(n10345) );
  CMPR32X1 U14032 ( .A(n10348), .B(n10347), .C(n10346), .CO(n10413), .S(n10419) );
  XNOR2XL U14033 ( .A(n9851), .B(n10341), .Y(n9655) );
  OAI22X1 U14034 ( .A0(n9963), .A1(n9665), .B0(n9631), .B1(n3180), .Y(n9658)
         );
  OAI22XL U14035 ( .A0(n10368), .A1(n9669), .B0(n9780), .B1(n9654), .Y(n9676)
         );
  ADDFX2 U14036 ( .A(n9884), .B(n9882), .CI(n9883), .CO(n9936), .S(n9935) );
  OAI22XL U14037 ( .A0(n9983), .A1(n9885), .B0(n9981), .B1(n9873), .Y(n9884)
         );
  CMPR32X1 U14038 ( .A(n9857), .B(n9856), .C(n9855), .CO(n10001), .S(n9858) );
  CMPR32X1 U14039 ( .A(n9969), .B(n9968), .C(n9967), .CO(n9993), .S(n10002) );
  OAI22XL U14040 ( .A0(n9966), .A1(n9834), .B0(n10159), .B1(n9965), .Y(n9968)
         );
  XNOR2X1 U14041 ( .A(n10324), .B(n9863), .Y(n9707) );
  XNOR2XL U14042 ( .A(n9851), .B(n10311), .Y(n9708) );
  NAND2BXL U14043 ( .AN(n9960), .B(M2_mult_x_15_n43), .Y(n9695) );
  NAND2BXL U14044 ( .AN(n9960), .B(n10339), .Y(n9737) );
  CMPR32X1 U14045 ( .A(n9822), .B(n9821), .C(n9820), .CO(n9809), .S(n10023) );
  XNOR2X1 U14046 ( .A(n9851), .B(n10387), .Y(n9630) );
  OAI22XL U14047 ( .A0(n10517), .A1(n6075), .B0(n9406), .B1(n10533), .Y(n9596)
         );
  INVXL U14048 ( .A(M2_b_17_), .Y(M2_U4_U1_or2_inv_0__14_) );
  NOR2XL U14049 ( .A(n5742), .B(M2_b_12_), .Y(M2_U4_U1_enc_tree_0__1__18_) );
  XNOR2XL U14050 ( .A(M2_a_17_), .B(n9863), .Y(n9419) );
  OAI22X1 U14051 ( .A0(n10368), .A1(n9252), .B0(n9780), .B1(n9265), .Y(n5245)
         );
  XNOR2X1 U14052 ( .A(M2_mult_x_15_n43), .B(n10311), .Y(n9297) );
  XNOR2X1 U14053 ( .A(n10339), .B(n10387), .Y(n9265) );
  AND2XL U14054 ( .A(n12311), .B(n12310), .Y(n12312) );
  NOR2BXL U14055 ( .AN(n3110), .B(n12119), .Y(n12149) );
  AND2X2 U14056 ( .A(n12118), .B(n4984), .Y(n12124) );
  OAI22XL U14057 ( .A0(n12595), .A1(n5516), .B0(n12597), .B1(n12009), .Y(
        n12016) );
  XNOR2XL U14058 ( .A(n12732), .B(n3110), .Y(n12003) );
  NAND2BXL U14059 ( .AN(n3110), .B(n12758), .Y(n11748) );
  OAI22XL U14060 ( .A0(n13838), .A1(n14198), .B0(n13781), .B1(n14208), .Y(
        n13857) );
  OR2X2 U14061 ( .A(n17881), .B(n18141), .Y(n5814) );
  OAI22XL U14062 ( .A0(n13156), .A1(n13899), .B0(n13058), .B1(n2997), .Y(
        n13162) );
  OAI22XL U14063 ( .A0(n13065), .A1(n13790), .B0(n13046), .B1(n13721), .Y(
        n13068) );
  ADDFX2 U14064 ( .A(n13091), .B(n4801), .CI(n13089), .CO(n13137), .S(n13136)
         );
  OAI22XL U14065 ( .A0(n13094), .A1(n2997), .B0(n13083), .B1(n13843), .Y(
        n13091) );
  OAI22XL U14066 ( .A0(n13155), .A1(n14044), .B0(n13171), .B1(n13974), .Y(
        n13178) );
  NOR2BXL U14067 ( .AN(n13049), .B(n14120), .Y(n13230) );
  OAI22XL U14068 ( .A0(n13284), .A1(n3173), .B0(n13224), .B1(n14080), .Y(
        n13263) );
  NAND2BXL U14069 ( .AN(n13049), .B(n14156), .Y(n13202) );
  OAI22XL U14070 ( .A0(n13208), .A1(n13721), .B0(n13170), .B1(n13790), .Y(
        n13210) );
  CMPR32X1 U14071 ( .A(n13217), .B(n13216), .C(n13215), .CO(n13274), .S(n13237) );
  OAI22XL U14072 ( .A0(n13208), .A1(n13790), .B0(n13218), .B1(n13721), .Y(
        n13216) );
  OAI22XL U14073 ( .A0(n13207), .A1(n14029), .B0(n13171), .B1(n14044), .Y(
        n13214) );
  OAI22XL U14074 ( .A0(n13267), .A1(n13899), .B0(n13220), .B1(n2997), .Y(
        n13290) );
  OAI22XL U14075 ( .A0(n13257), .A1(n13972), .B0(n13221), .B1(n13971), .Y(
        n13270) );
  OAI22XL U14076 ( .A0(n13315), .A1(n13721), .B0(n13285), .B1(n13790), .Y(
        n13330) );
  OAI22XL U14077 ( .A0(n13318), .A1(n3173), .B0(n13283), .B1(n14080), .Y(
        n13311) );
  OAI22XL U14078 ( .A0(n13317), .A1(n14120), .B0(n13279), .B1(n14121), .Y(
        n13325) );
  OAI22XL U14079 ( .A0(n13316), .A1(n14208), .B0(n13363), .B1(n14198), .Y(
        n13375) );
  NOR2BXL U14080 ( .AN(n13049), .B(n14227), .Y(n13374) );
  XNOR2XL U14081 ( .A(n14118), .B(n14030), .Y(n13421) );
  NAND2BXL U14082 ( .AN(n13049), .B(n14228), .Y(n13362) );
  XNOR2XL U14083 ( .A(n14235), .B(n13693), .Y(n13399) );
  NOR2BXL U14084 ( .AN(n13049), .B(n14268), .Y(n13433) );
  OAI22XL U14085 ( .A0(n13477), .A1(n13899), .B0(n13446), .B1(n2997), .Y(
        n13492) );
  NAND2XL U14086 ( .A(in_valid_d), .B(w1[134]), .Y(n11512) );
  INVXL U14087 ( .A(n25865), .Y(n13897) );
  XNOR2XL U14088 ( .A(n14306), .B(n14030), .Y(n13934) );
  XNOR2XL U14089 ( .A(n14235), .B(n25862), .Y(n13914) );
  XNOR2XL U14090 ( .A(n14265), .B(n14156), .Y(n13916) );
  OAI22XL U14091 ( .A0(n2993), .A1(n4565), .B0(n14356), .B1(n4567), .Y(n14026)
         );
  XNOR2X1 U14092 ( .A(n14265), .B(n25862), .Y(n14016) );
  CMPR32X1 U14093 ( .A(n14098), .B(n14097), .C(n14096), .CO(n14099), .S(n14166) );
  OAI22XL U14094 ( .A0(n14057), .A1(n14080), .B0(n3173), .B1(n25861), .Y(
        n14098) );
  OAI22XL U14095 ( .A0(n14135), .A1(n14268), .B0(n14079), .B1(n14282), .Y(
        n14125) );
  XOR2XL U14096 ( .A(n25884), .B(n3198), .Y(n4997) );
  OAI22XL U14097 ( .A0(n12352), .A1(n11892), .B0(n12222), .B1(n12233), .Y(
        n11912) );
  NOR2X1 U14098 ( .A(n15940), .B(n26004), .Y(n5047) );
  NOR2X1 U14099 ( .A(n15941), .B(n25901), .Y(n5048) );
  NOR2X1 U14100 ( .A(n15941), .B(n25905), .Y(n6088) );
  INVXL U14101 ( .A(n11485), .Y(n11486) );
  XNOR2X1 U14102 ( .A(n3199), .B(n12561), .Y(n16001) );
  XOR2X1 U14103 ( .A(n16614), .B(n5718), .Y(n15998) );
  OAI22X1 U14104 ( .A0(n18624), .A1(n17900), .B0(n18625), .B1(n17899), .Y(
        n17945) );
  OAI21X1 U14105 ( .A0(n18111), .A1(n5820), .B0(n5819), .Y(n17948) );
  XOR2X1 U14106 ( .A(n17908), .B(n4882), .Y(n17947) );
  ADDFX2 U14107 ( .A(n18148), .B(n4799), .CI(n18146), .CO(n18200), .S(n18199)
         );
  OAI22XL U14108 ( .A0(n18242), .A1(n18149), .B0(n18168), .B1(n18138), .Y(
        n18148) );
  OAI22XL U14109 ( .A0(n18242), .A1(n18178), .B0(n18168), .B1(n18149), .Y(
        n18189) );
  OAI22XL U14110 ( .A0(n18242), .A1(n18179), .B0(n18168), .B1(n18178), .Y(
        n18190) );
  NOR2BXL U14111 ( .AN(n2978), .B(n18238), .Y(n18192) );
  OAI22XL U14112 ( .A0(n18177), .A1(n18176), .B0(n18175), .B1(n18223), .Y(
        n18191) );
  AOI21XL U14113 ( .A0(n18174), .A1(n18170), .B0(n18173), .Y(n18186) );
  AND2XL U14114 ( .A(n18172), .B(n18171), .Y(n18173) );
  OAI22XL U14115 ( .A0(n5918), .A1(n18239), .B0(n18238), .B1(n18237), .Y(
        n18247) );
  OAI22XL U14116 ( .A0(n18107), .A1(n18236), .B0(n18235), .B1(n18234), .Y(
        n18248) );
  OAI22XL U14117 ( .A0(n5918), .A1(n18238), .B0(n18239), .B1(n18104), .Y(
        n18228) );
  OAI22X1 U14118 ( .A0(n18111), .A1(n18103), .B0(n18504), .B1(n6096), .Y(
        n18229) );
  OAI22X1 U14119 ( .A0(n18504), .A1(n5820), .B0(n17967), .B1(n18111), .Y(
        n17978) );
  OAI22XL U14120 ( .A0(n18111), .A1(n17999), .B0(n18504), .B1(n17967), .Y(
        n18004) );
  CMPR32X1 U14121 ( .A(n18019), .B(n18018), .C(n18017), .CO(n18016), .S(n18056) );
  OAI22XL U14122 ( .A0(n18541), .A1(n6129), .B0(n17995), .B1(n18539), .Y(
        n18023) );
  OAI22XL U14123 ( .A0(n18111), .A1(n18026), .B0(n18504), .B1(n17999), .Y(
        n18031) );
  NAND2BXL U14124 ( .AN(n2978), .B(n18453), .Y(n18008) );
  XNOR2X1 U14125 ( .A(n18500), .B(n18611), .Y(n5020) );
  NOR2BXL U14126 ( .AN(n13049), .B(n14298), .Y(n13515) );
  OAI22XL U14127 ( .A0(n13676), .A1(n14044), .B0(n13699), .B1(n13974), .Y(
        n13683) );
  XNOR2XL U14128 ( .A(n14027), .B(n25863), .Y(n13737) );
  XNOR2XL U14129 ( .A(n14357), .B(n4848), .Y(n13776) );
  NAND2XL U14130 ( .A(in_valid_d), .B(w1[129]), .Y(n13039) );
  OAI22XL U14131 ( .A0(n13714), .A1(n14080), .B0(n13793), .B1(n3173), .Y(
        n13772) );
  OAI22XL U14132 ( .A0(n13839), .A1(n14227), .B0(n13766), .B1(n14249), .Y(
        n13867) );
  OAI22XL U14133 ( .A0(n13841), .A1(n14080), .B0(n13874), .B1(n3173), .Y(
        n13877) );
  OAI22XL U14134 ( .A0(n13838), .A1(n14208), .B0(n13875), .B1(n14198), .Y(
        n13889) );
  INVXL U14135 ( .A(n8477), .Y(n8497) );
  INVXL U14136 ( .A(n19627), .Y(n19522) );
  NOR2X1 U14137 ( .A(n24092), .B(n19352), .Y(n19358) );
  AOI2BB2XL U14138 ( .B0(n3036), .B1(n19727), .A0N(n3036), .A1N(n19728), .Y(
        n19687) );
  OAI22XL U14139 ( .A0(n8510), .A1(n3017), .B0(n3040), .B1(n8509), .Y(n8621)
         );
  OAI22XL U14140 ( .A0(n8460), .A1(n3017), .B0(n3040), .B1(n8459), .Y(n8628)
         );
  OAI22XL U14141 ( .A0(n8475), .A1(n3017), .B0(n3040), .B1(n8474), .Y(n8632)
         );
  OAI22XL U14142 ( .A0(n8444), .A1(n3017), .B0(n3040), .B1(n8443), .Y(n8626)
         );
  INVXL U14143 ( .A(n8234), .Y(n8675) );
  INVXL U14144 ( .A(n8236), .Y(n8682) );
  INVXL U14145 ( .A(n8255), .Y(n8350) );
  INVXL U14146 ( .A(n8306), .Y(n8713) );
  NOR2XL U14147 ( .A(n8447), .B(n8513), .Y(n8515) );
  OAI22XL U14148 ( .A0(n8402), .A1(n3017), .B0(n3040), .B1(n8401), .Y(n8640)
         );
  OAI21XL U14149 ( .A0(n3160), .A1(n8325), .B0(n8324), .Y(n8647) );
  AOI21XL U14150 ( .A0(n8325), .A1(n8823), .B0(n3155), .Y(n8324) );
  OAI211XL U14151 ( .A0(n3154), .A1(n8489), .B0(n8295), .C0(n8323), .Y(n8325)
         );
  NAND2XL U14152 ( .A(n8476), .B(n3154), .Y(n8323) );
  OAI22XL U14153 ( .A0(n8327), .A1(n3017), .B0(n3040), .B1(n8326), .Y(n8646)
         );
  INVXL U14154 ( .A(n19366), .Y(n19811) );
  INVXL U14155 ( .A(n19554), .Y(n19584) );
  AOI2BB2XL U14156 ( .B0(n19727), .B1(n19542), .A0N(n19542), .A1N(n19726), .Y(
        n19790) );
  INVXL U14157 ( .A(n19385), .Y(n19480) );
  INVXL U14158 ( .A(n19370), .Y(n19816) );
  INVXL U14159 ( .A(n19364), .Y(n19803) );
  INVXL U14160 ( .A(n19435), .Y(n19842) );
  OAI21XL U14161 ( .A0(n3165), .A1(n19531), .B0(n19530), .Y(n19769) );
  AOI21XL U14162 ( .A0(n19531), .A1(n19952), .B0(n3164), .Y(n19530) );
  OAI21XL U14163 ( .A0(n19529), .A1(n19528), .B0(n19580), .Y(n19531) );
  OAI22XL U14164 ( .A0(n19533), .A1(n3100), .B0(n3041), .B1(n19532), .Y(n19768) );
  AOI21XL U14165 ( .A0(n19608), .A1(n3159), .B0(n19730), .Y(n19504) );
  NAND2XL U14166 ( .A(n19601), .B(n19807), .Y(n19503) );
  INVXL U14167 ( .A(n19484), .Y(n19509) );
  NAND2XL U14168 ( .A(n19546), .B(n19747), .Y(n19547) );
  NAND2XL U14169 ( .A(n19544), .B(n2996), .Y(n19545) );
  AOI22XL U14170 ( .A0(n19588), .A1(n4622), .B0(n19543), .B1(n19542), .Y(
        n19544) );
  INVXL U14171 ( .A(n19537), .Y(n19552) );
  OAI22XL U14172 ( .A0(n19599), .A1(n3100), .B0(n3041), .B1(n19598), .Y(n19703) );
  OAI22XL U14173 ( .A0(n19721), .A1(n3100), .B0(n19564), .B1(n19720), .Y(
        n19754) );
  OAI22XL U14174 ( .A0(n19737), .A1(n3100), .B0(n3041), .B1(n19736), .Y(n19756) );
  OAI22XL U14175 ( .A0(n19753), .A1(n3100), .B0(n19564), .B1(n19752), .Y(
        n19760) );
  INVXL U14176 ( .A(n19427), .Y(n19933) );
  OAI22XL U14177 ( .A0(n19456), .A1(n3100), .B0(n3041), .B1(n19455), .Y(n19774) );
  NOR2XL U14178 ( .A(n23208), .B(n23207), .Y(n19341) );
  AOI2BB2XL U14179 ( .B0(n3041), .B1(n19367), .A0N(n3041), .A1N(n19811), .Y(
        n19646) );
  NAND2XL U14180 ( .A(n3041), .B(n19393), .Y(n19394) );
  NAND2XL U14181 ( .A(n19564), .B(n19374), .Y(n19375) );
  NAND2XL U14182 ( .A(n2996), .B(n19640), .Y(n19651) );
  INVXL U14183 ( .A(n19616), .Y(n19650) );
  AOI2BB2XL U14184 ( .B0(n3041), .B1(n19436), .A0N(n3041), .A1N(n19842), .Y(
        n19676) );
  AOI2BB2XL U14185 ( .B0(n3041), .B1(n19365), .A0N(n3041), .A1N(n19803), .Y(
        n19659) );
  NAND2XL U14186 ( .A(n3041), .B(n19390), .Y(n19391) );
  AOI2BB2XL U14187 ( .B0(n3041), .B1(n19561), .A0N(n3041), .A1N(n19721), .Y(
        n19616) );
  NAND2XL U14188 ( .A(n19564), .B(n19438), .Y(n19439) );
  AOI2BB2XL U14189 ( .B0(n3041), .B1(n19568), .A0N(n3041), .A1N(n19753), .Y(
        n19632) );
  AOI2BB2XL U14190 ( .B0(n3041), .B1(n19384), .A0N(n3041), .A1N(n19456), .Y(
        n19627) );
  NOR2XL U14191 ( .A(n3167), .B(n15264), .Y(n15266) );
  INVXL U14192 ( .A(n14997), .Y(n15098) );
  INVXL U14193 ( .A(n15005), .Y(n15414) );
  INVXL U14194 ( .A(n15416), .Y(n15417) );
  OAI22XL U14195 ( .A0(n15210), .A1(n3156), .B0(n3016), .B1(n15209), .Y(n15419) );
  INVXL U14196 ( .A(n14980), .Y(n15423) );
  AOI2BB2XL U14197 ( .B0(n15558), .B1(n14983), .A0N(n15190), .A1N(n15431), .Y(
        n15320) );
  AOI2BB2XL U14198 ( .B0(n15190), .B1(n14981), .A0N(n15190), .A1N(n15423), .Y(
        n15338) );
  AOI2BB2XL U14199 ( .B0(n15190), .B1(n15057), .A0N(n15190), .A1N(n15462), .Y(
        n15334) );
  NOR2X1 U14200 ( .A(n3090), .B(n3016), .Y(n15336) );
  NAND2XL U14201 ( .A(n15190), .B(n15066), .Y(n15067) );
  NAND2XL U14202 ( .A(n15190), .B(n15059), .Y(n15060) );
  NAND2XL U14203 ( .A(n15190), .B(n15103), .Y(n15104) );
  NAND2XL U14204 ( .A(n15190), .B(n15172), .Y(n15173) );
  NAND2XL U14205 ( .A(n15190), .B(n15002), .Y(n15003) );
  NAND2XL U14206 ( .A(n15190), .B(n15177), .Y(n15178) );
  AOI2BB2XL U14207 ( .B0(n15558), .B1(n14996), .A0N(n15558), .A1N(n15076), .Y(
        n15288) );
  NAND2XL U14208 ( .A(n15190), .B(n15106), .Y(n15107) );
  INVXL U14209 ( .A(n21958), .Y(n21652) );
  INVXL U14210 ( .A(n21558), .Y(n21559) );
  INVXL U14211 ( .A(n21898), .Y(n21635) );
  OAI22XL U14212 ( .A0(n15260), .A1(n3101), .B0(n15190), .B1(n15259), .Y(
        n15368) );
  OAI22XL U14213 ( .A0(n15207), .A1(n3101), .B0(n15558), .B1(n15206), .Y(
        n15375) );
  OAI21XL U14214 ( .A0(n14967), .A1(n15149), .B0(n15148), .Y(n15388) );
  OAI21XL U14215 ( .A0(n15147), .A1(n15146), .B0(n15256), .Y(n15149) );
  AOI21XL U14216 ( .A0(n3090), .A1(n15349), .B0(n15145), .Y(n15146) );
  OAI22XL U14217 ( .A0(n15151), .A1(n3101), .B0(n15558), .B1(n15150), .Y(
        n15387) );
  INVXL U14218 ( .A(n15225), .Y(n15243) );
  INVXL U14219 ( .A(n15142), .Y(n15143) );
  AOI21XL U14220 ( .A0(n15268), .A1(n15313), .B0(n15355), .Y(n15122) );
  NAND2XL U14221 ( .A(n15263), .B(n3090), .Y(n15121) );
  INVXL U14222 ( .A(n15102), .Y(n15127) );
  NAND2XL U14223 ( .A(n15162), .B(n15313), .Y(n15163) );
  AOI22XL U14224 ( .A0(n15248), .A1(n6194), .B0(n15160), .B1(n3016), .Y(n15162) );
  INVXL U14225 ( .A(n15159), .Y(n15160) );
  INVXL U14226 ( .A(n15549), .Y(n15165) );
  INVXL U14227 ( .A(n15154), .Y(n15170) );
  INVXL U14228 ( .A(n14982), .Y(n15431) );
  INVXL U14229 ( .A(n15065), .Y(n15543) );
  INVXL U14230 ( .A(n15062), .Y(n15538) );
  INVXL U14231 ( .A(n15058), .Y(n15522) );
  INVXL U14232 ( .A(n14986), .Y(n15436) );
  OAI22XL U14233 ( .A0(n15076), .A1(n3101), .B0(n15008), .B1(n15075), .Y(
        n15393) );
  NAND2XL U14234 ( .A(n21659), .B(n3171), .Y(n21573) );
  NAND2XL U14235 ( .A(n21609), .B(n3037), .Y(n21610) );
  AOI22XL U14236 ( .A0(n21646), .A1(n3172), .B0(n21608), .B1(n3096), .Y(n21609) );
  INVXL U14237 ( .A(n21607), .Y(n21608) );
  INVXL U14238 ( .A(n21989), .Y(n21612) );
  OAI22XL U14239 ( .A0(n21791), .A1(n3042), .B0(n3020), .B1(n21200), .Y(n21813) );
  OAI22XL U14240 ( .A0(n21810), .A1(n3042), .B0(n23116), .B1(n21201), .Y(
        n21817) );
  AOI2BB2XL U14241 ( .B0(n3172), .B1(n21767), .A0N(n3172), .A1N(n21766), .Y(
        n21840) );
  NAND2XL U14242 ( .A(n21778), .B(n3096), .Y(n21747) );
  OAI21XL U14243 ( .A0(n21854), .A1(n21599), .B0(n21598), .Y(n21826) );
  AOI21XL U14244 ( .A0(n21599), .A1(n3222), .B0(n21849), .Y(n21598) );
  AOI22XL U14245 ( .A0(n21803), .A1(n22011), .B0(n21596), .B1(n21595), .Y(
        n21597) );
  OAI22XL U14246 ( .A0(n21601), .A1(n3042), .B0(n3020), .B1(n21224), .Y(n21825) );
  OAI22XL U14247 ( .A0(n21531), .A1(n3042), .B0(n3020), .B1(n21225), .Y(n21831) );
  INVXL U14248 ( .A(n21855), .Y(n21856) );
  OAI22XL U14249 ( .A0(n8379), .A1(n3017), .B0(n3040), .B1(n8378), .Y(n8638)
         );
  OAI22XL U14250 ( .A0(n8421), .A1(n3017), .B0(n3040), .B1(n8420), .Y(n8636)
         );
  NAND2XL U14251 ( .A(n6217), .B(y10[18]), .Y(n8046) );
  XNOR2X1 U14252 ( .A(M3_mult_x_15_a_17_), .B(n5430), .Y(n11649) );
  XNOR2XL U14253 ( .A(n12282), .B(n3202), .Y(n11652) );
  INVXL U14254 ( .A(n12282), .Y(n12285) );
  XNOR2X1 U14255 ( .A(n12758), .B(n3197), .Y(n11782) );
  AOI21XL U14256 ( .A0(n23021), .A1(n11071), .B0(n22887), .Y(n22580) );
  ADDFX2 U14257 ( .A(n7574), .B(n7573), .CI(n7572), .CO(n7578), .S(n7557) );
  OAI22XL U14258 ( .A0(n4592), .A1(n7555), .B0(n3046), .B1(n25869), .Y(n7573)
         );
  NOR2XL U14259 ( .A(n11073), .B(n3219), .Y(n22555) );
  INVXL U14260 ( .A(n22567), .Y(n22554) );
  INVXL U14261 ( .A(n22553), .Y(n22568) );
  NAND2XL U14262 ( .A(n11073), .B(n3219), .Y(n22556) );
  AOI21XL U14263 ( .A0(n22927), .A1(n3218), .B0(n21073), .Y(n21074) );
  OAI2BB1XL U14264 ( .A0N(n11071), .A1N(n22700), .B0(n22701), .Y(n21073) );
  CMPR32X1 U14265 ( .A(n7631), .B(n7630), .C(n7629), .CO(n7649), .S(n7637) );
  INVXL U14266 ( .A(n25876), .Y(n7631) );
  OAI22XL U14267 ( .A0(n7633), .A1(n23221), .B0(n7634), .B1(n7615), .Y(n7630)
         );
  ADDFX2 U14268 ( .A(n7592), .B(n7591), .CI(n7590), .CO(n7612), .S(n7579) );
  INVXL U14269 ( .A(n7621), .Y(n7592) );
  OAI22XL U14270 ( .A0(n7633), .A1(n7570), .B0(n7589), .B1(n6300), .Y(n7591)
         );
  OAI21XL U14271 ( .A0(n5124), .A1(n7588), .B0(n5106), .Y(n7618) );
  CMPR32X1 U14272 ( .A(n7586), .B(n7585), .C(n7584), .CO(n7624), .S(n7583) );
  XOR2XL U14273 ( .A(n3054), .B(n11214), .Y(n10759) );
  XNOR2XL U14274 ( .A(n3053), .B(n11213), .Y(n10760) );
  XNOR2XL U14275 ( .A(n11214), .B(n11213), .Y(n10758) );
  AOI222XL U14276 ( .A0(n22892), .A1(n11058), .B0(n22708), .B1(n23151), .C0(
        n22891), .C1(n10789), .Y(n22882) );
  INVXL U14277 ( .A(n22931), .Y(n22911) );
  XOR2XL U14278 ( .A(n3055), .B(n21078), .Y(n21081) );
  XNOR2XL U14279 ( .A(n3054), .B(n21079), .Y(n21082) );
  XNOR2XL U14280 ( .A(n21079), .B(n21078), .Y(n21080) );
  AOI222XL U14281 ( .A0(n23003), .A1(n11074), .B0(n22969), .B1(n3219), .C0(
        n23001), .C1(n11073), .Y(n22669) );
  INVXL U14282 ( .A(n22870), .Y(n22871) );
  AOI222XL U14283 ( .A0(n23152), .A1(n3220), .B0(n23093), .B1(n22867), .C0(
        n23150), .C1(n10775), .Y(n22868) );
  AOI222XL U14284 ( .A0(n22892), .A1(n11059), .B0(n22708), .B1(n11058), .C0(
        n22891), .C1(n23151), .Y(n22884) );
  AOI222XL U14285 ( .A0(n23152), .A1(n10789), .B0(n23093), .B1(n3220), .C0(
        n23150), .C1(n26496), .Y(n23147) );
  AOI21XL U14286 ( .A0(n23021), .A1(n3218), .B0(n22888), .Y(n22889) );
  OAI2BB1XL U14287 ( .A0N(n11071), .A1N(n22887), .B0(n22886), .Y(n22888) );
  AOI222XL U14288 ( .A0(n23003), .A1(n23109), .B0(n22969), .B1(n11062), .C0(
        n23001), .C1(n3217), .Y(n22964) );
  AOI222XL U14289 ( .A0(n22928), .A1(n23151), .B0(n22700), .B1(n10789), .C0(
        n22927), .C1(n3220), .Y(n22878) );
  AOI222XL U14290 ( .A0(n22892), .A1(n26496), .B0(n22708), .B1(n10775), .C0(
        n22891), .C1(n10769), .Y(n22876) );
  INVXL U14291 ( .A(n23001), .Y(n22599) );
  INVXL U14292 ( .A(n22976), .Y(n22539) );
  NAND2XL U14293 ( .A(n11074), .B(n3219), .Y(n22526) );
  XNOR2XL U14294 ( .A(n21059), .B(n21058), .Y(n21070) );
  AOI21XL U14295 ( .A0(n22976), .A1(n11071), .B0(n22980), .Y(n21065) );
  AOI21XL U14296 ( .A0(n22976), .A1(n3218), .B0(n22564), .Y(n22565) );
  OAI2BB1XL U14297 ( .A0N(n11071), .A1N(n22980), .B0(n22981), .Y(n22564) );
  OAI22XL U14298 ( .A0(n4592), .A1(n7531), .B0(n3046), .B1(n7555), .Y(n7552)
         );
  CMPR32X1 U14299 ( .A(n7473), .B(n7472), .C(n7471), .CO(n7496), .S(n7469) );
  XOR2XL U14300 ( .A(n22796), .B(n3221), .Y(M6_mult_x_15_n1203) );
  XOR2XL U14301 ( .A(n22815), .B(n3053), .Y(M6_mult_x_15_n1178) );
  XOR2XL U14302 ( .A(n22955), .B(n3221), .Y(M6_mult_x_15_n1202) );
  XOR2XL U14303 ( .A(n22821), .B(n3221), .Y(M6_mult_x_15_n1200) );
  AOI222XL U14304 ( .A0(n22988), .A1(n10789), .B0(n22980), .B1(n3220), .C0(
        n22976), .C1(n26496), .Y(n22808) );
  NAND2XL U14305 ( .A(n9109), .B(n3218), .Y(n22507) );
  INVXL U14306 ( .A(n22941), .Y(n22942) );
  OAI2BB2XL U14307 ( .B0(n23073), .B1(n3225), .A0N(n22987), .A1N(n23093), .Y(
        n22941) );
  INVXL U14308 ( .A(n10812), .Y(n10814) );
  XNOR2XL U14309 ( .A(n10872), .B(n10871), .Y(n22869) );
  NAND2XL U14310 ( .A(n10870), .B(n11049), .Y(n10871) );
  INVXL U14311 ( .A(n11047), .Y(n10870) );
  XNOR2XL U14312 ( .A(n22780), .B(n22779), .Y(n23135) );
  NAND2XL U14313 ( .A(n22778), .B(n22777), .Y(n22779) );
  AOI21XL U14314 ( .A0(n22775), .A1(n22774), .B0(n22773), .Y(n22780) );
  INVXL U14315 ( .A(n22776), .Y(n22778) );
  NOR2XL U14316 ( .A(n11141), .B(n11143), .Y(n22500) );
  NOR2XL U14317 ( .A(n11144), .B(n11146), .Y(n22553) );
  NOR2XL U14318 ( .A(n11152), .B(n11154), .Y(n22605) );
  NOR2XL U14319 ( .A(n11166), .B(n11168), .Y(n11131) );
  NAND2XL U14320 ( .A(n7329), .B(M0_U4_U1_enc_tree_3__3__24_), .Y(n7332) );
  INVXL U14321 ( .A(M0_U4_U1_enc_tree_3__3__16_), .Y(n7329) );
  ADDFX2 U14322 ( .A(n6696), .B(n6695), .CI(n6694), .CO(n6465), .S(n6711) );
  AND2XL U14323 ( .A(n6590), .B(n6589), .Y(n6594) );
  AND2XL U14324 ( .A(n6592), .B(n6591), .Y(n6593) );
  ADDFX2 U14325 ( .A(n6654), .B(n6653), .CI(n6652), .CO(n6661), .S(n6660) );
  XOR3X2 U14326 ( .A(n6509), .B(n6508), .C(n6507), .Y(n6667) );
  OAI21XL U14327 ( .A0(n6508), .A1(n6509), .B0(n6507), .Y(n5629) );
  OAI22XL U14328 ( .A0(n6540), .A1(n7460), .B0(n7535), .B1(n6539), .Y(n6683)
         );
  INVXL U14329 ( .A(n6533), .Y(n5575) );
  OAI22XL U14330 ( .A0(n7535), .A1(n6312), .B0(n6311), .B1(n7556), .Y(n6339)
         );
  OAI21X1 U14331 ( .A0(n6346), .A1(n7695), .B0(n5123), .Y(n6351) );
  OR2X2 U14332 ( .A(n6780), .B(n7093), .Y(n5130) );
  XNOR2XL U14333 ( .A(n3209), .B(n25875), .Y(n5131) );
  NAND2BXL U14334 ( .AN(n6944), .B(n23219), .Y(n6747) );
  XNOR2X1 U14335 ( .A(n7534), .B(M0_a_12_), .Y(n5572) );
  XNOR2XL U14336 ( .A(n25866), .B(n25873), .Y(n6835) );
  XOR2X1 U14337 ( .A(n6028), .B(n7615), .Y(n6027) );
  NAND2XL U14338 ( .A(n12945), .B(M3_U3_U1_enc_tree_3__3__24_), .Y(n12946) );
  INVXL U14339 ( .A(M3_U3_U1_enc_tree_3__3__16_), .Y(n12945) );
  INVXL U14340 ( .A(M3_U3_U1_enc_tree_1__2__12_), .Y(
        M3_U3_U1_enc_tree_1__3__8_) );
  OR2XL U14341 ( .A(M3_U3_U1_or2_tree_1__2__16_), .B(
        M3_U3_U1_or2_tree_1__2__24_), .Y(n26151) );
  AND2XL U14342 ( .A(M3_U3_U1_enc_tree_1__1__12_), .B(
        M3_U3_U1_enc_tree_1__1__14_), .Y(n25990) );
  OR2XL U14343 ( .A(M3_U3_U1_enc_tree_2__2__16_), .B(
        M3_U3_U1_enc_tree_2__2__24_), .Y(n26203) );
  AOI21XL U14344 ( .A0(n4875), .A1(data[37]), .B0(n4963), .Y(n4962) );
  AOI21XL U14345 ( .A0(n12225), .A1(M3_a_10_), .B0(n5970), .Y(
        M3_U3_U1_enc_tree_0__1__22_) );
  XNOR2X1 U14346 ( .A(n18638), .B(n5430), .Y(n17500) );
  XNOR2X1 U14347 ( .A(n18468), .B(n12561), .Y(n17508) );
  XOR2XL U14348 ( .A(n3053), .B(n11217), .Y(n10784) );
  XNOR2XL U14349 ( .A(n11217), .B(n11219), .Y(n10783) );
  AOI222XL U14350 ( .A0(n23023), .A1(n3219), .B0(n22887), .B1(n11073), .C0(
        n23021), .C1(n11063), .Y(n22851) );
  AOI222XL U14351 ( .A0(n22932), .A1(n3218), .B0(n22904), .B1(n23089), .C0(
        n22931), .C1(n11074), .Y(n22730) );
  XOR2XL U14352 ( .A(n22856), .B(n3056), .Y(M6_mult_x_15_n1096) );
  XNOR2XL U14353 ( .A(n22643), .B(n21087), .Y(n23155) );
  NAND2XL U14354 ( .A(n21086), .B(n22641), .Y(n21087) );
  INVXL U14355 ( .A(n22642), .Y(n21086) );
  AOI222XL U14356 ( .A0(n22988), .A1(n23109), .B0(n22980), .B1(n11062), .C0(
        n22976), .C1(n3217), .Y(n22849) );
  INVXL U14357 ( .A(n22925), .Y(n22926) );
  AOI222XL U14358 ( .A0(n23152), .A1(n26496), .B0(n23093), .B1(n10775), .C0(
        n23150), .C1(n10769), .Y(n22923) );
  AOI222XL U14359 ( .A0(n23003), .A1(n3219), .B0(n22969), .B1(n11073), .C0(
        n23001), .C1(n11063), .Y(n22919) );
  AOI222XL U14360 ( .A0(n23023), .A1(n3218), .B0(n22887), .B1(n23089), .C0(
        n23021), .C1(n11074), .Y(n22734) );
  AOI21XL U14361 ( .A0(n22931), .A1(n11071), .B0(n22904), .Y(n22783) );
  XOR2XL U14362 ( .A(n22930), .B(n3058), .Y(M6_mult_x_15_n1069) );
  AOI222XL U14363 ( .A0(n23023), .A1(n11074), .B0(n22887), .B1(n3219), .C0(
        n23021), .C1(n11073), .Y(n22789) );
  AOI222XL U14364 ( .A0(n22928), .A1(n11058), .B0(n22700), .B1(n23151), .C0(
        n22927), .C1(n10789), .Y(n22787) );
  AOI222XL U14365 ( .A0(n22988), .A1(n3217), .B0(n22980), .B1(n23022), .C0(
        n22976), .C1(n11059), .Y(n22841) );
  INVXL U14366 ( .A(n22952), .Y(n22833) );
  AOI222XL U14367 ( .A0(n22892), .A1(n10789), .B0(n22708), .B1(n3220), .C0(
        n22891), .C1(n26496), .Y(n22755) );
  INVXL U14368 ( .A(n22827), .Y(n22828) );
  AOI222XL U14369 ( .A0(n23152), .A1(n10775), .B0(n23093), .B1(n10769), .C0(
        n23150), .C1(n23002), .Y(n22826) );
  AND2XL U14370 ( .A(n16656), .B(n16655), .Y(n16657) );
  XNOR2X1 U14371 ( .A(n5858), .B(n5546), .Y(n16485) );
  ADDFX2 U14372 ( .A(n16389), .B(n16388), .CI(n16387), .CO(n16394), .S(n16456)
         );
  OAI22XL U14373 ( .A0(n16942), .A1(n16353), .B0(n16688), .B1(n16359), .Y(
        n16388) );
  OAI22XL U14374 ( .A0(n3102), .A1(n16352), .B0(n16332), .B1(n16351), .Y(
        n16389) );
  OAI22X1 U14375 ( .A0(n17060), .A1(n16349), .B0(n17061), .B1(n5704), .Y(
        n16385) );
  NAND2X1 U14376 ( .A(n5857), .B(n5856), .Y(n16406) );
  XOR2X1 U14377 ( .A(n3199), .B(n16965), .Y(n16117) );
  XNOR2X1 U14378 ( .A(n3199), .B(M3_mult_x_15_b_9_), .Y(n16048) );
  OAI22X1 U14379 ( .A0(n17060), .A1(n5706), .B0(n17061), .B1(n16102), .Y(
        n16442) );
  CMPR32X1 U14380 ( .A(n16420), .B(n16419), .C(n16418), .CO(n16820), .S(n16449) );
  OAI22X1 U14381 ( .A0(n17074), .A1(n16072), .B0(n16375), .B1(n5693), .Y(
        n16110) );
  OAI22X1 U14382 ( .A0(n17074), .A1(n5693), .B0(n16375), .B1(n16007), .Y(
        n16093) );
  INVXL U14383 ( .A(M5_U3_U1_enc_tree_1__2__12_), .Y(
        M5_U3_U1_enc_tree_1__3__8_) );
  OR2XL U14384 ( .A(M5_U3_U1_or2_tree_1__2__16_), .B(
        M5_U3_U1_or2_tree_1__2__24_), .Y(n26206) );
  AND2XL U14385 ( .A(M5_U3_U1_enc_tree_1__1__12_), .B(
        M5_U3_U1_enc_tree_1__1__14_), .Y(n25982) );
  OR2XL U14386 ( .A(M5_U3_U1_enc_tree_2__2__16_), .B(
        M5_U3_U1_enc_tree_2__2__24_), .Y(n26196) );
  NOR2X1 U14387 ( .A(n15942), .B(n6181), .Y(n5435) );
  INVXL U14388 ( .A(M4_U3_U1_enc_tree_2__2__24_), .Y(M4_U3_U1_or2_inv_2__24_)
         );
  NOR2XL U14389 ( .A(M4_a_19_), .B(M4_a_18_), .Y(M4_U3_U1_enc_tree_1__1__12_)
         );
  NOR2XL U14390 ( .A(n11074), .B(n9109), .Y(n22530) );
  INVXL U14391 ( .A(n22526), .Y(n22527) );
  INVXL U14392 ( .A(n22500), .Y(n22528) );
  NAND2XL U14393 ( .A(n11074), .B(n9109), .Y(n22531) );
  NAND2XL U14394 ( .A(n10794), .B(n10793), .Y(n11222) );
  NAND2XL U14395 ( .A(w2[32]), .B(n23973), .Y(n10794) );
  NAND2XL U14396 ( .A(w2[64]), .B(valid[0]), .Y(n10793) );
  NAND2XL U14397 ( .A(n10755), .B(n10754), .Y(n11213) );
  NAND2XL U14398 ( .A(w2[70]), .B(valid[0]), .Y(n10754) );
  NAND2XL U14399 ( .A(w2[38]), .B(n23973), .Y(n10755) );
  NAND2XL U14400 ( .A(n10757), .B(n10756), .Y(n11214) );
  NAND2XL U14401 ( .A(w2[71]), .B(valid[0]), .Y(n10756) );
  NAND2XL U14402 ( .A(w2[39]), .B(n23973), .Y(n10757) );
  NAND2XL U14403 ( .A(n11196), .B(n11195), .Y(n21078) );
  NAND2XL U14404 ( .A(w2[74]), .B(valid[0]), .Y(n11195) );
  NAND2XL U14405 ( .A(w2[42]), .B(n23973), .Y(n11196) );
  AOI2BB1XL U14406 ( .A0N(n11186), .A1N(n21058), .B0(n22990), .Y(n11192) );
  NAND2XL U14407 ( .A(n11199), .B(n11198), .Y(n21079) );
  NAND2XL U14408 ( .A(w2[73]), .B(valid[0]), .Y(n11198) );
  NAND2XL U14409 ( .A(w2[41]), .B(n23973), .Y(n11199) );
  NAND2XL U14410 ( .A(n10782), .B(n10781), .Y(n11217) );
  NAND2XL U14411 ( .A(w2[36]), .B(n23973), .Y(n10782) );
  NAND2XL U14412 ( .A(w2[68]), .B(valid[0]), .Y(n10781) );
  NAND3XL U14413 ( .A(n26195), .B(y11[2]), .C(n23973), .Y(n10747) );
  AOI2BB1XL U14414 ( .A0N(n11157), .A1N(n11156), .B0(n11155), .Y(n11158) );
  AOI2BB1XL U14415 ( .A0N(n11154), .A1N(n11153), .B0(n11152), .Y(n11156) );
  AOI2BB1XL U14416 ( .A0N(n11151), .A1N(n11150), .B0(n23022), .Y(n11153) );
  AOI2BB1XL U14417 ( .A0N(n11149), .A1N(n11148), .B0(n11147), .Y(n11150) );
  NAND2XL U14418 ( .A(w2[51]), .B(n3501), .Y(n11172) );
  NAND2XL U14419 ( .A(w2[83]), .B(valid[0]), .Y(n11171) );
  NAND2XL U14420 ( .A(w2[82]), .B(valid[0]), .Y(n11173) );
  NAND2XL U14421 ( .A(w2[50]), .B(n3501), .Y(n11174) );
  XNOR2XL U14422 ( .A(n22492), .B(n22491), .Y(n22493) );
  NAND2XL U14423 ( .A(n22496), .B(n11076), .Y(n22505) );
  NAND2XL U14424 ( .A(w2[85]), .B(valid[0]), .Y(n11085) );
  NAND2XL U14425 ( .A(w2[53]), .B(n23973), .Y(n11086) );
  NAND2XL U14426 ( .A(w2[86]), .B(valid[0]), .Y(n11087) );
  NAND2XL U14427 ( .A(w2[54]), .B(n23973), .Y(n11088) );
  XNOR2XL U14428 ( .A(n16614), .B(n3202), .Y(n16125) );
  INVXL U14429 ( .A(n5642), .Y(n5640) );
  XNOR2X1 U14430 ( .A(n3203), .B(n3048), .Y(n16253) );
  CMPR32X1 U14431 ( .A(n16222), .B(n16221), .C(n16220), .CO(n16232), .S(n16213) );
  OAI22X1 U14432 ( .A0(n17148), .A1(n3108), .B0(n17147), .B1(n3049), .Y(n16206) );
  OAI22X1 U14433 ( .A0(n16164), .A1(n17060), .B0(n17061), .B1(n16201), .Y(
        n16209) );
  XOR2XL U14434 ( .A(n3201), .B(n16909), .Y(n5329) );
  NOR2XL U14435 ( .A(n8610), .B(n3157), .Y(n8538) );
  NAND2XL U14436 ( .A(n3040), .B(n8264), .Y(n8265) );
  NAND2XL U14437 ( .A(n8482), .B(n8244), .Y(n8245) );
  NAND2XL U14438 ( .A(n8161), .B(n8408), .Y(n8409) );
  NAND2XL U14439 ( .A(n8482), .B(n8241), .Y(n8242) );
  INVXL U14440 ( .A(n8572), .Y(n8578) );
  INVXL U14441 ( .A(n8526), .Y(n8573) );
  NAND2XL U14442 ( .A(n8482), .B(n8261), .Y(n8262) );
  NAND2XL U14443 ( .A(n8482), .B(n8309), .Y(n8310) );
  OAI21XL U14444 ( .A0(n8482), .A1(n8794), .B0(n8317), .Y(n8534) );
  NAND2XL U14445 ( .A(n8482), .B(n8316), .Y(n8317) );
  NAND2XL U14446 ( .A(n8482), .B(n8425), .Y(n8426) );
  INVXL U14447 ( .A(n19441), .Y(n19918) );
  INVXL U14448 ( .A(n19444), .Y(n19923) );
  INVXL U14449 ( .A(n19425), .Y(n19928) );
  CMPR32X1 U14450 ( .A(n7478), .B(n7477), .C(n7476), .CO(n7494), .S(n7457) );
  CMPR32X1 U14451 ( .A(n7296), .B(n7295), .C(n7294), .CO(n7458), .S(n7276) );
  CMPR32X1 U14452 ( .A(n10307), .B(n10306), .C(n10305), .CO(n10433), .S(n10302) );
  NAND2XL U14453 ( .A(n5543), .B(n10171), .Y(n5539) );
  NAND2XL U14454 ( .A(n5304), .B(n9478), .Y(n5299) );
  CMPR32X1 U14455 ( .A(n9541), .B(n9540), .C(n9539), .CO(n9567), .S(n9530) );
  OAI22XL U14456 ( .A0(n10541), .A1(n9536), .B0(n10329), .B1(n9580), .Y(n9572)
         );
  OAI22XL U14457 ( .A0(n9966), .A1(n9501), .B0(n10159), .B1(n9550), .Y(n9535)
         );
  OAI2BB1XL U14458 ( .A0N(n10369), .A1N(n10368), .B0(n10339), .Y(n10389) );
  OAI22XL U14459 ( .A0(n9504), .A1(n10381), .B0(n10496), .B1(n10404), .Y(
        n10398) );
  INVXL U14460 ( .A(n10335), .Y(n9103) );
  OAI22XL U14461 ( .A0(n9504), .A1(n4808), .B0(n10496), .B1(n5202), .Y(n10491)
         );
  INVXL U14462 ( .A(n15047), .Y(n15548) );
  INVXL U14463 ( .A(n15052), .Y(n15559) );
  NAND2X1 U14464 ( .A(n5144), .B(n5143), .Y(n9692) );
  NAND2XL U14465 ( .A(n9677), .B(n5148), .Y(n5143) );
  NAND2XL U14466 ( .A(n5145), .B(n9676), .Y(n5144) );
  NAND2BXL U14467 ( .AN(n9677), .B(n5146), .Y(n5145) );
  AND2XL U14468 ( .A(n9931), .B(n9930), .Y(n9932) );
  NAND2XL U14469 ( .A(n9797), .B(n5188), .Y(n5184) );
  NAND2BXL U14470 ( .AN(n9797), .B(n5186), .Y(n5185) );
  OAI22XL U14471 ( .A0(n9966), .A1(n9817), .B0(n10159), .B1(n9798), .Y(n10019)
         );
  NOR2BXL U14472 ( .AN(n9960), .B(n10659), .Y(n9327) );
  OAI22XL U14473 ( .A0(n10541), .A1(n9396), .B0(n10329), .B1(n9302), .Y(n9325)
         );
  OAI22X1 U14474 ( .A0(n10296), .A1(n9600), .B0(n9959), .B1(n9433), .Y(n9623)
         );
  OAI22XL U14475 ( .A0(n9590), .A1(n9589), .B0(n9877), .B1(n9439), .Y(n9626)
         );
  CMPR32X1 U14476 ( .A(n9606), .B(n9605), .C(n9604), .CO(n10089), .S(n10077)
         );
  OAI22XL U14477 ( .A0(n9966), .A1(n9612), .B0(n10159), .B1(n9443), .Y(n9606)
         );
  CMPR32X1 U14478 ( .A(n9449), .B(n9448), .C(n9447), .CO(n9430), .S(n10088) );
  OAI22X1 U14479 ( .A0(n10368), .A1(n9446), .B0(n9780), .B1(n9382), .Y(n9449)
         );
  OAI22XL U14480 ( .A0(n9445), .A1(n9444), .B0(n9906), .B1(n9384), .Y(n9448)
         );
  OAI22X1 U14481 ( .A0(n9433), .A1(n10296), .B0(n9959), .B1(n5376), .Y(n9452)
         );
  OR2XL U14482 ( .A(M2_U4_U1_enc_tree_2__2__16_), .B(
        M2_U4_U1_enc_tree_2__2__24_), .Y(n26197) );
  OR2XL U14483 ( .A(M2_U3_U1_enc_tree_2__2__16_), .B(
        M2_U3_U1_enc_tree_2__2__24_), .Y(n26204) );
  NAND2XL U14484 ( .A(n9285), .B(n9284), .Y(n5349) );
  ADDFX2 U14485 ( .A(n9401), .B(n9400), .CI(n9399), .CO(n9428), .S(n10072) );
  OAI22X1 U14486 ( .A0(n9321), .A1(n9959), .B0(n10296), .B1(n5376), .Y(n9400)
         );
  OAI22XL U14487 ( .A0(n9551), .A1(n9421), .B0(n9838), .B1(n9320), .Y(n9401)
         );
  NAND2BXL U14488 ( .AN(n9423), .B(n5533), .Y(n5532) );
  OAI22XL U14489 ( .A0(n11878), .A1(n12633), .B0(n12635), .B1(n6040), .Y(
        n11894) );
  XNOR2XL U14490 ( .A(n12233), .B(n12803), .Y(n11763) );
  XOR2XL U14491 ( .A(n12233), .B(n6112), .Y(n11636) );
  XNOR2X1 U14492 ( .A(n12732), .B(M3_mult_x_15_b_9_), .Y(n11783) );
  OAI22X1 U14493 ( .A0(n12635), .A1(n11688), .B0(n12513), .B1(n11687), .Y(
        n11702) );
  INVXL U14494 ( .A(n12352), .Y(n5326) );
  OAI22X1 U14495 ( .A0(n12717), .A1(n11722), .B0(n12718), .B1(n11649), .Y(
        n5964) );
  XOR2XL U14496 ( .A(n25884), .B(n6112), .Y(n12534) );
  OAI21XL U14497 ( .A0(n12386), .A1(n12387), .B0(n12385), .Y(n5791) );
  CMPR32X1 U14498 ( .A(n12140), .B(n12139), .C(n12138), .CO(n12133), .S(n12215) );
  XNOR2X1 U14499 ( .A(n12519), .B(n3190), .Y(n11670) );
  XNOR2X1 U14500 ( .A(n3204), .B(n12561), .Y(n11850) );
  OAI22XL U14501 ( .A0(n12635), .A1(n11852), .B0(n12513), .B1(n11792), .Y(
        n11854) );
  OAI22X1 U14502 ( .A0(n12717), .A1(n12004), .B0(n12718), .B1(n11843), .Y(
        n12047) );
  OAI22XL U14503 ( .A0(n11994), .A1(n12352), .B0(n12222), .B1(n6105), .Y(
        n12050) );
  XNOR2XL U14504 ( .A(n12282), .B(M3_mult_x_15_b_19_), .Y(n11794) );
  XOR2XL U14505 ( .A(n12282), .B(n6112), .Y(n11793) );
  XNOR2XL U14506 ( .A(n25884), .B(n3049), .Y(n11844) );
  OAI22X1 U14507 ( .A0(n12715), .A1(n12002), .B0(n12525), .B1(n6115), .Y(
        n11998) );
  NOR2BXL U14508 ( .AN(n3110), .B(n12760), .Y(n12000) );
  OAI21X2 U14509 ( .A0(n25911), .A1(n15942), .B0(n5419), .Y(M3_a_16_) );
  NOR2X1 U14510 ( .A(n17167), .B(n26017), .Y(n5958) );
  XNOR2X1 U14511 ( .A(n12751), .B(n5997), .Y(n12575) );
  NOR2X1 U14512 ( .A(n4860), .B(n25916), .Y(n4920) );
  OAI21XL U14513 ( .A0(n26011), .A1(n15940), .B0(n4930), .Y(n4929) );
  NOR2X1 U14514 ( .A(n4860), .B(n25914), .Y(n4946) );
  NAND2XL U14515 ( .A(n11479), .B(data[51]), .Y(n4930) );
  NAND2XL U14516 ( .A(n18083), .B(n18429), .Y(n5463) );
  OAI22XL U14517 ( .A0(n14075), .A1(n14208), .B0(n14089), .B1(n14198), .Y(
        n14087) );
  OAI22XL U14518 ( .A0(n14071), .A1(n6191), .B0(n14078), .B1(n14298), .Y(
        n14083) );
  OAI22XL U14519 ( .A0(n14069), .A1(n14282), .B0(n14079), .B1(n14251), .Y(
        n14084) );
  OAI22X1 U14520 ( .A0(n14157), .A1(n5510), .B0(n14120), .B1(n14156), .Y(
        n14132) );
  CMPR32X1 U14521 ( .A(n18507), .B(n18506), .C(n18505), .CO(n18493), .S(n18529) );
  OAI22XL U14522 ( .A0(n18659), .A1(n18542), .B0(n17832), .B1(n18431), .Y(
        n18506) );
  OAI22XL U14523 ( .A0(n18083), .A1(n17879), .B0(n4649), .B1(n18429), .Y(
        n17885) );
  XNOR2X1 U14524 ( .A(n18118), .B(n3201), .Y(n17581) );
  XNOR2XL U14525 ( .A(n18500), .B(M3_mult_x_15_b_13_), .Y(n17539) );
  XNOR2X1 U14526 ( .A(n18503), .B(n3198), .Y(n17538) );
  OAI22XL U14527 ( .A0(n18541), .A1(n17862), .B0(n5769), .B1(n18539), .Y(
        n17876) );
  OAI22XL U14528 ( .A0(n18111), .A1(n17892), .B0(n18504), .B1(n17717), .Y(
        n17878) );
  OAI22X2 U14529 ( .A0(n18652), .A1(n17873), .B0(n17872), .B1(n17871), .Y(
        n17890) );
  OAI22X1 U14530 ( .A0(n18652), .A1(n17871), .B0(n17872), .B1(n17681), .Y(
        n17867) );
  AND2XL U14531 ( .A(n13131), .B(n13130), .Y(n13132) );
  ADDFX2 U14532 ( .A(n13426), .B(n13425), .CI(n13424), .CO(n13501), .S(n13452)
         );
  OAI22XL U14533 ( .A0(n13364), .A1(n14044), .B0(n13421), .B1(n13974), .Y(
        n13426) );
  CMPR32X1 U14534 ( .A(n13527), .B(n13526), .C(n13525), .CO(n13571), .S(n13516) );
  CMPR32X1 U14535 ( .A(n13530), .B(n13529), .C(n13528), .CO(n13570), .S(n13519) );
  CMPR32X1 U14536 ( .A(n13472), .B(n13471), .C(n13470), .CO(n13546), .S(n13487) );
  OAI22XL U14537 ( .A0(n13493), .A1(n13972), .B0(n13451), .B1(n13971), .Y(
        n13470) );
  OAI22XL U14538 ( .A0(n13482), .A1(n13721), .B0(n13450), .B1(n13790), .Y(
        n13471) );
  XNOR2XL U14539 ( .A(n14265), .B(n4848), .Y(n13565) );
  XNOR2XL U14540 ( .A(n14028), .B(n25862), .Y(n13541) );
  XNOR2XL U14541 ( .A(n14027), .B(n25862), .Y(n13566) );
  OAI22XL U14542 ( .A0(n13493), .A1(n13971), .B0(n13506), .B1(n13972), .Y(
        n13537) );
  NAND2X1 U14543 ( .A(n3123), .B(w1[150]), .Y(n11547) );
  NAND2XL U14544 ( .A(n14365), .B(M1_U3_U1_enc_tree_3__3__24_), .Y(n14368) );
  INVXL U14545 ( .A(M1_U3_U1_enc_tree_3__3__16_), .Y(n14365) );
  OR2XL U14546 ( .A(M1_U3_U1_or2_tree_1__2__16_), .B(
        M1_U3_U1_or2_tree_1__2__24_), .Y(n26210) );
  INVXL U14547 ( .A(M1_U3_U1_enc_tree_1__2__12_), .Y(
        M1_U3_U1_enc_tree_1__3__8_) );
  INVXL U14548 ( .A(M1_U4_U1_enc_tree_1__2__12_), .Y(
        M1_U4_U1_enc_tree_1__3__8_) );
  OR2XL U14549 ( .A(M1_U4_U1_or2_tree_1__2__16_), .B(
        M1_U4_U1_or2_tree_1__2__24_), .Y(n26211) );
  AND2XL U14550 ( .A(M1_U4_U1_enc_tree_1__1__12_), .B(
        M1_U4_U1_enc_tree_1__1__14_), .Y(n25983) );
  OR2XL U14551 ( .A(M1_U4_U1_enc_tree_2__2__16_), .B(
        M1_U4_U1_enc_tree_2__2__24_), .Y(n26202) );
  AND2XL U14552 ( .A(M1_U3_U1_enc_tree_1__1__12_), .B(
        M1_U3_U1_enc_tree_1__1__14_), .Y(n25987) );
  OR2XL U14553 ( .A(M1_U3_U1_enc_tree_2__2__16_), .B(
        M1_U3_U1_enc_tree_2__2__24_), .Y(n26199) );
  XOR2X1 U14554 ( .A(M3_mult_x_15_n1682), .B(n18658), .Y(n5455) );
  XNOR2XL U14555 ( .A(n18468), .B(M3_mult_x_15_b_13_), .Y(n17636) );
  XNOR2X1 U14556 ( .A(n18604), .B(n3190), .Y(n17619) );
  CMPR32X1 U14557 ( .A(n17838), .B(n17837), .C(n17836), .CO(n18526), .S(n17839) );
  OAI22XL U14558 ( .A0(n18111), .A1(n17791), .B0(n18504), .B1(n18503), .Y(
        n17837) );
  OAI22X1 U14559 ( .A0(n18721), .A1(n3197), .B0(n17512), .B1(
        M3_mult_x_15_n1682), .Y(n17786) );
  CMPR32X1 U14560 ( .A(n17755), .B(n17754), .C(n17753), .CO(n17773), .S(n17803) );
  NAND2XL U14561 ( .A(n13928), .B(n13927), .Y(n4874) );
  OAI22XL U14562 ( .A0(n13917), .A1(n14282), .B0(n13973), .B1(n14251), .Y(
        n13966) );
  OAI2BB1X1 U14563 ( .A0N(n14056), .A1N(n14055), .B0(n5490), .Y(n14171) );
  OAI21XL U14564 ( .A0(n14055), .A1(n14056), .B0(n14054), .Y(n5490) );
  OAI22XL U14565 ( .A0(n14190), .A1(n14227), .B0(n14159), .B1(n14249), .Y(
        n14199) );
  CMPR32X1 U14566 ( .A(n14155), .B(n14154), .C(n14153), .CO(n14183), .S(n14139) );
  OAI22XL U14567 ( .A0(n14135), .A1(n14282), .B0(n14158), .B1(n14251), .Y(
        n14153) );
  OAI22XL U14568 ( .A0(n14134), .A1(n14208), .B0(n14148), .B1(n14198), .Y(
        n14154) );
  INVXL U14569 ( .A(n4997), .Y(n4995) );
  XNOR2X1 U14570 ( .A(n3204), .B(n3202), .Y(n11958) );
  OAI21XL U14571 ( .A0(n12715), .A1(n11918), .B0(n4907), .Y(n11954) );
  NOR2XL U14572 ( .A(n3205), .B(n16475), .Y(n15980) );
  OAI21X1 U14573 ( .A0(n15966), .A1(n17060), .B0(n5641), .Y(n15988) );
  NAND2BXL U14574 ( .AN(n18076), .B(n6128), .Y(n6127) );
  INVXL U14575 ( .A(n18077), .Y(n6128) );
  CMPR32X1 U14576 ( .A(n17701), .B(n17700), .C(n17699), .CO(n17704), .S(n18338) );
  OAI22X1 U14577 ( .A0(n18522), .A1(n17678), .B0(n3195), .B1(n17600), .Y(
        n17701) );
  OAI22XL U14578 ( .A0(n18721), .A1(M3_mult_x_15_b_3_), .B0(n17512), .B1(
        n11499), .Y(n17559) );
  OAI22XL U14579 ( .A0(n17551), .A1(n5893), .B0(n17552), .B1(n18541), .Y(
        n17564) );
  OAI22XL U14580 ( .A0(M3_mult_x_15_b_1_), .A1(n17512), .B0(n2978), .B1(n18721), .Y(n17541) );
  OAI22X1 U14581 ( .A0(n17539), .A1(n18083), .B0(n18429), .B1(n5020), .Y(
        n17550) );
  INVXL U14582 ( .A(n14236), .Y(n14217) );
  OAI22XL U14583 ( .A0(n14208), .A1(n25862), .B0(n14198), .B1(n14197), .Y(
        n14215) );
  OAI22XL U14584 ( .A0(n2993), .A1(n14235), .B0(n14289), .B1(n14266), .Y(
        n14216) );
  INVXL U14585 ( .A(n14266), .Y(n14248) );
  OAI22XL U14586 ( .A0(n14249), .A1(n14228), .B0(n14227), .B1(n3019), .Y(
        n14246) );
  OAI22XL U14587 ( .A0(n2993), .A1(n14265), .B0(n14289), .B1(n25864), .Y(
        n14247) );
  OAI22XL U14588 ( .A0(n14233), .A1(n14268), .B0(n14210), .B1(n14282), .Y(
        n14229) );
  OAI22XL U14589 ( .A0(n14190), .A1(n14249), .B0(n14214), .B1(n14250), .Y(
        n14211) );
  OAI22XL U14590 ( .A0(n14188), .A1(n14282), .B0(n14210), .B1(n14251), .Y(
        n14213) );
  OAI22XL U14591 ( .A0(n13576), .A1(n14120), .B0(n13539), .B1(n14121), .Y(
        n13573) );
  XNOR3X2 U14592 ( .A(n5215), .B(n13730), .C(n13731), .Y(n13711) );
  NAND2XL U14593 ( .A(n13731), .B(n5214), .Y(n5212) );
  OAI22XL U14594 ( .A0(n14263), .A1(n14291), .B0(n14253), .B1(n6191), .Y(
        n14260) );
  OAI22XL U14595 ( .A0(n14263), .A1(n6191), .B0(n14283), .B1(n14298), .Y(
        n14281) );
  OAI2BB1XL U14596 ( .A0N(n14268), .A1N(n14282), .B0(n25863), .Y(n14294) );
  OAI22XL U14597 ( .A0(n14283), .A1(n6191), .B0(n14298), .B1(n23173), .Y(
        n14293) );
  OAI22XL U14598 ( .A0(n8497), .A1(n3017), .B0(n3040), .B1(n8496), .Y(n8619)
         );
  INVXL U14599 ( .A(n8621), .Y(n4815) );
  NAND2XL U14600 ( .A(n8633), .B(n8632), .Y(n8893) );
  OAI22XL U14601 ( .A0(n8675), .A1(n3017), .B0(n3040), .B1(n8674), .Y(n8697)
         );
  AOI21XL U14602 ( .A0(n8680), .A1(n8823), .B0(n3155), .Y(n8679) );
  OAI211XL U14603 ( .A0(n3154), .A1(n8678), .B0(n8295), .C0(n8677), .Y(n8680)
         );
  OAI22XL U14604 ( .A0(n8682), .A1(n3017), .B0(n3040), .B1(n8681), .Y(n8699)
         );
  AOI21XL U14605 ( .A0(n8690), .A1(n8823), .B0(n3155), .Y(n8689) );
  NAND2XL U14606 ( .A(n8295), .B(n8688), .Y(n8690) );
  OAI22XL U14607 ( .A0(n8692), .A1(n3017), .B0(n3040), .B1(n8691), .Y(n8705)
         );
  OAI22XL U14608 ( .A0(n8350), .A1(n3017), .B0(n3040), .B1(n8349), .Y(n8648)
         );
  OAI22XL U14609 ( .A0(n8713), .A1(n3017), .B0(n3040), .B1(n8712), .Y(n8714)
         );
  INVXL U14610 ( .A(n8308), .Y(n8773) );
  INVXL U14611 ( .A(n8315), .Y(n8794) );
  INVXL U14612 ( .A(n8312), .Y(n8789) );
  INVXL U14613 ( .A(n8296), .Y(n8799) );
  INVXL U14614 ( .A(n8298), .Y(n8804) );
  OAI21XL U14615 ( .A0(n3160), .A1(n8658), .B0(n8657), .Y(n8694) );
  AOI21XL U14616 ( .A0(n8658), .A1(n8823), .B0(n3155), .Y(n8657) );
  NAND2XL U14617 ( .A(n8295), .B(n8656), .Y(n8658) );
  AOI22XL U14618 ( .A0(n8655), .A1(n3086), .B0(n8654), .B1(n3154), .Y(n8656)
         );
  OAI22XL U14619 ( .A0(n8660), .A1(n3017), .B0(n3040), .B1(n8659), .Y(n8693)
         );
  AOI21XL U14620 ( .A0(n8665), .A1(n8823), .B0(n3155), .Y(n8664) );
  NAND2XL U14621 ( .A(n8295), .B(n8663), .Y(n8665) );
  AOI22XL U14622 ( .A0(n8662), .A1(n3086), .B0(n8661), .B1(n3154), .Y(n8663)
         );
  OAI22XL U14623 ( .A0(n8667), .A1(n3017), .B0(n3040), .B1(n8666), .Y(n8695)
         );
  NAND2XL U14624 ( .A(n8295), .B(n8683), .Y(n8685) );
  OAI22XL U14625 ( .A0(n8687), .A1(n3017), .B0(n3040), .B1(n8686), .Y(n8703)
         );
  NOR2XL U14626 ( .A(n8924), .B(n8927), .Y(n8929) );
  INVXL U14627 ( .A(n8931), .Y(n8642) );
  INVXL U14628 ( .A(n8925), .Y(n8643) );
  OAI22XL U14629 ( .A0(n19811), .A1(n3100), .B0(n3041), .B1(n19810), .Y(n19828) );
  OAI22XL U14630 ( .A0(n19821), .A1(n3100), .B0(n3041), .B1(n19820), .Y(n19834) );
  OAI22XL U14631 ( .A0(n19584), .A1(n3100), .B0(n3041), .B1(n19583), .Y(n19701) );
  OAI22XL U14632 ( .A0(n19795), .A1(n3100), .B0(n3041), .B1(n19794), .Y(n19824) );
  AOI21XL U14633 ( .A0(n19478), .A1(n19952), .B0(n3164), .Y(n19477) );
  NAND2XL U14634 ( .A(n19424), .B(n19476), .Y(n19478) );
  AOI22XL U14635 ( .A0(n19591), .A1(n3159), .B0(n19592), .B1(n19807), .Y(
        n19476) );
  OAI22XL U14636 ( .A0(n19480), .A1(n3100), .B0(n3041), .B1(n19479), .Y(n19776) );
  OAI22XL U14637 ( .A0(n19788), .A1(n3100), .B0(n3041), .B1(n19787), .Y(n19822) );
  OAI22XL U14638 ( .A0(n19816), .A1(n3100), .B0(n3041), .B1(n19815), .Y(n19832) );
  OAI22XL U14639 ( .A0(n19803), .A1(n3100), .B0(n3041), .B1(n19802), .Y(n19826) );
  OAI22XL U14640 ( .A0(n19902), .A1(n3100), .B0(n3041), .B1(n19901), .Y(n19904) );
  OAI22XL U14641 ( .A0(n19842), .A1(n3100), .B0(n3041), .B1(n19841), .Y(n19843) );
  NAND2XL U14642 ( .A(n19769), .B(n19768), .Y(n20060) );
  NOR2XL U14643 ( .A(n20053), .B(n20056), .Y(n20058) );
  OAI22XL U14644 ( .A0(n19509), .A1(n3100), .B0(n3041), .B1(n19508), .Y(n19766) );
  OAI22XL U14645 ( .A0(n19552), .A1(n3100), .B0(n3041), .B1(n19551), .Y(n19764) );
  INVXL U14646 ( .A(n19431), .Y(n19938) );
  INVX1 U14647 ( .A(n19432), .Y(n19937) );
  NAND4BXL U14648 ( .AN(n19674), .B(n19673), .C(n19672), .D(n19671), .Y(n19680) );
  AOI21XL U14649 ( .A0(n2996), .A1(n3094), .B0(n19623), .Y(n19626) );
  OAI22XL U14650 ( .A0(n15098), .A1(n3101), .B0(n15008), .B1(n15097), .Y(
        n15395) );
  NAND2XL U14651 ( .A(n15046), .B(n15403), .Y(n15405) );
  AOI22XL U14652 ( .A0(n15402), .A1(n3034), .B0(n15401), .B1(n3090), .Y(n15403) );
  OAI22XL U14653 ( .A0(n15407), .A1(n3101), .B0(n15558), .B1(n15406), .Y(
        n15442) );
  NAND2XL U14654 ( .A(n15046), .B(n15410), .Y(n15412) );
  AOI22XL U14655 ( .A0(n15409), .A1(n3034), .B0(n15408), .B1(n3090), .Y(n15410) );
  OAI22XL U14656 ( .A0(n15414), .A1(n3101), .B0(n15008), .B1(n15413), .Y(
        n15444) );
  OAI22XL U14657 ( .A0(n15423), .A1(n3101), .B0(n15008), .B1(n15422), .Y(
        n15446) );
  INVXL U14658 ( .A(n15049), .Y(n15553) );
  OAI22XL U14659 ( .A0(n21657), .A1(n3042), .B0(n3020), .B1(n21194), .Y(n21758) );
  NAND2XL U14660 ( .A(n21840), .B(n3171), .Y(n21770) );
  OAI22XL U14661 ( .A0(n21640), .A1(n3042), .B0(n3020), .B1(n21193), .Y(n21756) );
  NOR2XL U14662 ( .A(n3095), .B(n21660), .Y(n21663) );
  NAND2XL U14663 ( .A(n21181), .B(n21180), .Y(n21656) );
  NAND2XL U14664 ( .A(n21192), .B(n21191), .Y(n21639) );
  INVXL U14665 ( .A(n21619), .Y(n21640) );
  INVXL U14666 ( .A(n23120), .Y(n21486) );
  INVXL U14667 ( .A(n21639), .Y(n21193) );
  INVXL U14668 ( .A(n21656), .Y(n21194) );
  NAND2XL U14669 ( .A(n21183), .B(n21182), .Y(n21620) );
  NAND3XL U14670 ( .A(cs[0]), .B(cs[1]), .C(target_temp[1]), .Y(n21182) );
  NAND2XL U14671 ( .A(n21188), .B(n21187), .Y(n21623) );
  NAND3XL U14672 ( .A(cs[0]), .B(cs[1]), .C(target_temp[2]), .Y(n21187) );
  INVXL U14673 ( .A(n21790), .Y(n21200) );
  NAND2XL U14674 ( .A(n21329), .B(temp0[6]), .Y(n21214) );
  NOR2XL U14675 ( .A(n15674), .B(n15677), .Y(n15679) );
  NAND2XL U14676 ( .A(n15388), .B(n15387), .Y(n15681) );
  OAI22XL U14677 ( .A0(n15243), .A1(n3101), .B0(n15558), .B1(n15242), .Y(
        n15366) );
  INVXL U14678 ( .A(n14967), .Y(n15415) );
  AOI2BB2XL U14679 ( .B0(n15354), .B1(n3016), .A0N(n15353), .A1N(n3016), .Y(
        n15356) );
  OAI22XL U14680 ( .A0(n15198), .A1(n6194), .B0(n3016), .B1(n15195), .Y(n15358) );
  OAI22XL U14681 ( .A0(n15127), .A1(n3101), .B0(n15190), .B1(n15126), .Y(
        n15385) );
  OAI22XL U14682 ( .A0(n15170), .A1(n3101), .B0(n15008), .B1(n15169), .Y(
        n15383) );
  OAI211XL U14683 ( .A0(n3090), .A1(n15427), .B0(n15046), .C0(n15426), .Y(
        n15429) );
  OAI22XL U14684 ( .A0(n15431), .A1(n3101), .B0(n15558), .B1(n15430), .Y(
        n15448) );
  OAI22XL U14685 ( .A0(n15543), .A1(n3101), .B0(n15558), .B1(n15542), .Y(
        n15562) );
  NAND2XL U14686 ( .A(n15046), .B(n15534), .Y(n15536) );
  NAND2XL U14687 ( .A(n15046), .B(n15518), .Y(n15520) );
  OAI22XL U14688 ( .A0(n15522), .A1(n3101), .B0(n15558), .B1(n15521), .Y(
        n15524) );
  NAND2XL U14689 ( .A(n15046), .B(n15432), .Y(n15434) );
  OAI22XL U14690 ( .A0(n15436), .A1(n3101), .B0(n15008), .B1(n15435), .Y(
        n15452) );
  INVXL U14691 ( .A(n14988), .Y(n15441) );
  INVXL U14692 ( .A(n15056), .Y(n15462) );
  OAI22XL U14693 ( .A0(n21579), .A1(n3042), .B0(n3020), .B1(n21220), .Y(n21823) );
  OAI22XL U14694 ( .A0(n21617), .A1(n3042), .B0(n3020), .B1(n21219), .Y(n21821) );
  OAI21XL U14695 ( .A0(n21854), .A1(n21551), .B0(n21550), .Y(n21834) );
  AOI21XL U14696 ( .A0(n21551), .A1(n3222), .B0(n21849), .Y(n21550) );
  OAI211XL U14697 ( .A0(n3171), .A1(n21650), .B0(n21506), .C0(n21549), .Y(
        n21551) );
  NAND2XL U14698 ( .A(n21641), .B(n3171), .Y(n21549) );
  OAI22XL U14699 ( .A0(n21553), .A1(n3042), .B0(n3020), .B1(n21260), .Y(n21833) );
  OAI21XL U14700 ( .A0(n21854), .A1(n21851), .B0(n21850), .Y(n21885) );
  NAND2XL U14701 ( .A(n21506), .B(n21848), .Y(n21851) );
  AOI22XL U14702 ( .A0(n21847), .A1(n4618), .B0(n21846), .B1(n3171), .Y(n21848) );
  OAI22XL U14703 ( .A0(n21853), .A1(n21429), .B0(n3020), .B1(n21265), .Y(
        n21884) );
  OAI21XL U14704 ( .A0(n21854), .A1(n21843), .B0(n21842), .Y(n21883) );
  AOI21XL U14705 ( .A0(n21843), .A1(n3222), .B0(n21849), .Y(n21842) );
  NAND2XL U14706 ( .A(n21506), .B(n21841), .Y(n21843) );
  AOI22XL U14707 ( .A0(n21840), .A1(n3037), .B0(n21839), .B1(n3171), .Y(n21841) );
  OAI22XL U14708 ( .A0(n21845), .A1(n3042), .B0(n3020), .B1(n21261), .Y(n21882) );
  OAI21XL U14709 ( .A0(n21854), .A1(n21874), .B0(n21873), .Y(n21893) );
  AOI21XL U14710 ( .A0(n21874), .A1(n3222), .B0(n21849), .Y(n21873) );
  NAND2XL U14711 ( .A(n21506), .B(n21872), .Y(n21874) );
  OAI22XL U14712 ( .A0(n21876), .A1(n3042), .B0(n3020), .B1(n21274), .Y(n21892) );
  INVXL U14713 ( .A(n21508), .Y(n21988) );
  NAND2X2 U14714 ( .A(n21723), .B(n21500), .Y(n21787) );
  INVX1 U14715 ( .A(n21673), .Y(n21500) );
  OAI21XL U14716 ( .A0(n21854), .A1(n21869), .B0(n21868), .Y(n21889) );
  AOI21XL U14717 ( .A0(n21869), .A1(n3222), .B0(n21849), .Y(n21868) );
  OAI211XL U14718 ( .A0(n3171), .A1(n21867), .B0(n21506), .C0(n21866), .Y(
        n21869) );
  OAI22XL U14719 ( .A0(n21871), .A1(n3042), .B0(n3020), .B1(n21273), .Y(n21888) );
  OAI21XL U14720 ( .A0(n21854), .A1(n21879), .B0(n21878), .Y(n21895) );
  AOI21XL U14721 ( .A0(n21879), .A1(n3222), .B0(n21849), .Y(n21878) );
  NAND2XL U14722 ( .A(n21506), .B(n21877), .Y(n21879) );
  OAI22XL U14723 ( .A0(n21881), .A1(n3042), .B0(n3020), .B1(n21278), .Y(n21894) );
  OAI21XL U14724 ( .A0(n21854), .A1(n21900), .B0(n21899), .Y(n21904) );
  AOI21XL U14725 ( .A0(n21900), .A1(n3222), .B0(n21849), .Y(n21899) );
  NAND2XL U14726 ( .A(n21506), .B(n21898), .Y(n21900) );
  OAI22XL U14727 ( .A0(n21902), .A1(n3042), .B0(n3020), .B1(n21279), .Y(n21903) );
  NOR2XL U14728 ( .A(n22111), .B(n22114), .Y(n22116) );
  NAND2XL U14729 ( .A(n21826), .B(n21825), .Y(n22118) );
  OAI22XL U14730 ( .A0(n21863), .A1(n3042), .B0(n3020), .B1(n21266), .Y(n21886) );
  NAND2XL U14731 ( .A(n8639), .B(n8638), .Y(n8925) );
  INVXL U14732 ( .A(n8924), .Y(n8915) );
  OAI22XL U14733 ( .A0(n17087), .A1(n17059), .B0(n16375), .B1(n17073), .Y(
        n17069) );
  OAI22XL U14734 ( .A0(n17092), .A1(n17071), .B0(n17099), .B1(n17086), .Y(
        n17085) );
  XOR2XL U14735 ( .A(n22628), .B(n3058), .Y(M6_mult_x_15_n1064) );
  INVXL U14736 ( .A(n23140), .Y(M6_mult_x_15_n1017) );
  XOR2XL U14737 ( .A(n22840), .B(n3055), .Y(M6_mult_x_15_n1112) );
  XOR2XL U14738 ( .A(n22813), .B(n3119), .Y(M6_mult_x_15_n1040) );
  NAND2XL U14739 ( .A(n16972), .B(n5672), .Y(n5668) );
  XOR2XL U14740 ( .A(n22676), .B(n3056), .Y(M6_mult_x_15_n1089) );
  XOR2XL U14741 ( .A(n22830), .B(n3054), .Y(M6_mult_x_15_n1137) );
  XOR2XL U14742 ( .A(n22748), .B(n3055), .Y(M6_mult_x_15_n1113) );
  XOR2XL U14743 ( .A(n22581), .B(n3054), .Y(M6_mult_x_15_n1138) );
  XOR2XL U14744 ( .A(n22754), .B(n3058), .Y(M6_mult_x_15_n1066) );
  INVXL U14745 ( .A(n23156), .Y(M6_mult_x_15_n1019) );
  XOR2XL U14746 ( .A(n22686), .B(n3055), .Y(M6_mult_x_15_n1114) );
  XOR2XL U14747 ( .A(n22786), .B(n3056), .Y(M6_mult_x_15_n1090) );
  XOR2XL U14748 ( .A(n22832), .B(n3119), .Y(M6_mult_x_15_n1042) );
  INVXL U14749 ( .A(n22578), .Y(n22579) );
  XOR2XL U14750 ( .A(n22656), .B(n3055), .Y(M6_mult_x_15_n1111) );
  XOR2XL U14751 ( .A(n22794), .B(n3058), .Y(M6_mult_x_15_n1063) );
  INVXL U14752 ( .A(n23146), .Y(M6_mult_x_15_n1016) );
  INVXL U14753 ( .A(n23105), .Y(M6_mult_x_15_n1011) );
  INVXL U14754 ( .A(n22927), .Y(n21060) );
  XOR2XL U14755 ( .A(n22542), .B(n3058), .Y(n22543) );
  AOI21XL U14756 ( .A0(n22927), .A1(n11071), .B0(n22700), .Y(n22541) );
  CMPR32X1 U14757 ( .A(n7643), .B(n7642), .C(n7641), .CO(n7688), .S(n7648) );
  OAI2BB1XL U14758 ( .A0N(n7634), .A1N(n7633), .B0(n6299), .Y(n7641) );
  OAI22XL U14759 ( .A0(n7829), .A1(n25875), .B0(n7828), .B1(n25874), .Y(n7643)
         );
  OAI2BB2XL U14760 ( .B0(n5124), .B1(n7632), .A0N(n5122), .A1N(n7644), .Y(
        n7642) );
  ADDFX2 U14761 ( .A(n7637), .B(n7636), .CI(n7635), .CO(n7638), .S(n7655) );
  ADDFX2 U14762 ( .A(n7614), .B(n7613), .CI(n7612), .CO(n7656), .S(n7622) );
  OAI22XL U14763 ( .A0(n7829), .A1(n25876), .B0(n7828), .B1(n7646), .Y(n7614)
         );
  ADDFX2 U14764 ( .A(n7624), .B(n7623), .CI(n7622), .CO(n7654), .S(n7651) );
  XOR2XL U14765 ( .A(n22540), .B(n3056), .Y(M6_mult_x_15_n1083) );
  INVXL U14766 ( .A(n23108), .Y(M6_mult_x_15_n1012) );
  ADDFX2 U14767 ( .A(n7595), .B(n7594), .CI(n7593), .CO(n7604), .S(n7607) );
  XOR2XL U14768 ( .A(n22782), .B(n3053), .Y(M6_mult_x_15_n1175) );
  AOI222XL U14769 ( .A0(n22932), .A1(n11063), .B0(n22904), .B1(n23109), .C0(
        n22931), .C1(n11062), .Y(n22695) );
  NOR2XL U14770 ( .A(M6_mult_x_15_n667), .B(M6_mult_x_15_n674), .Y(n10921) );
  XOR2XL U14771 ( .A(n3221), .B(n11221), .Y(n10799) );
  XNOR2XL U14772 ( .A(n11222), .B(n11221), .Y(n10798) );
  AOI222XL U14773 ( .A0(n23023), .A1(n23109), .B0(n22887), .B1(n11062), .C0(
        n23021), .C1(n3217), .Y(n22859) );
  AOI222XL U14774 ( .A0(n22932), .A1(n3219), .B0(n22904), .B1(n11073), .C0(
        n22931), .C1(n11063), .Y(n22901) );
  XOR2XL U14775 ( .A(n22717), .B(n22716), .Y(n22728) );
  AOI222XL U14776 ( .A0(n22928), .A1(n10775), .B0(n22700), .B1(n10769), .C0(
        n22927), .C1(n23002), .Y(n22715) );
  AOI222XL U14777 ( .A0(n23003), .A1(n11059), .B0(n22969), .B1(n11058), .C0(
        n23001), .C1(n23151), .Y(n22611) );
  AOI222XL U14778 ( .A0(n23003), .A1(n3217), .B0(n22969), .B1(n23022), .C0(
        n23001), .C1(n11059), .Y(n22804) );
  AOI222XL U14779 ( .A0(n22932), .A1(n11074), .B0(n22904), .B1(n3219), .C0(
        n22931), .C1(n11073), .Y(n22770) );
  NAND2XL U14780 ( .A(w2[75]), .B(valid[0]), .Y(n11193) );
  NAND2XL U14781 ( .A(w2[43]), .B(n23973), .Y(n11194) );
  XOR2XL U14782 ( .A(n22895), .B(n3119), .Y(M6_mult_x_15_n1051) );
  XOR2XL U14783 ( .A(n21077), .B(n22716), .Y(M6_mult_x_15_n1075) );
  INVXL U14784 ( .A(n22940), .Y(n22949) );
  AOI222XL U14785 ( .A0(n23152), .A1(n10749), .B0(n23093), .B1(n3116), .C0(
        n23150), .C1(n22987), .Y(n22939) );
  AND2XL U14786 ( .A(M0_U3_U1_enc_tree_1__1__12_), .B(
        M0_U3_U1_enc_tree_1__1__14_), .Y(n25986) );
  OR2XL U14787 ( .A(M0_U3_U1_enc_tree_2__2__16_), .B(
        M0_U3_U1_enc_tree_2__2__24_), .Y(n26201) );
  AND2XL U14788 ( .A(M0_U4_U1_enc_tree_1__1__12_), .B(
        M0_U4_U1_enc_tree_1__1__14_), .Y(n25988) );
  OR2XL U14789 ( .A(M0_U4_U1_enc_tree_2__2__16_), .B(
        M0_U4_U1_enc_tree_2__2__24_), .Y(n26198) );
  INVXL U14790 ( .A(M0_U3_U1_enc_tree_3__3__16_), .Y(n7330) );
  INVXL U14791 ( .A(n7332), .Y(n7335) );
  INVXL U14792 ( .A(M0_U4_U1_enc_tree_1__2__12_), .Y(
        M0_U4_U1_enc_tree_1__3__8_) );
  OR2XL U14793 ( .A(M0_U4_U1_or2_tree_1__2__16_), .B(
        M0_U4_U1_or2_tree_1__2__24_), .Y(n26148) );
  OR2XL U14794 ( .A(M0_U3_U1_or2_tree_1__2__16_), .B(
        M0_U3_U1_or2_tree_1__2__24_), .Y(n26147) );
  INVXL U14795 ( .A(M0_U3_U1_enc_tree_1__2__12_), .Y(
        M0_U3_U1_enc_tree_1__3__8_) );
  INVXL U14796 ( .A(M0_U3_U1_enc_tree_2__4__16_), .Y(n7352) );
  INVXL U14797 ( .A(M0_U4_U1_enc_tree_2__4__16_), .Y(n7353) );
  AOI22XL U14798 ( .A0(n7337), .A1(n7333), .B0(n7335), .B1(n7334), .Y(n7339)
         );
  NAND2XL U14799 ( .A(n7332), .B(n7331), .Y(n7333) );
  INVXL U14800 ( .A(n7334), .Y(n7331) );
  NOR2XL U14801 ( .A(n7341), .B(n7342), .Y(n7340) );
  INVXL U14802 ( .A(M0_U4_U1_enc_tree_1__4__16_), .Y(n7349) );
  INVXL U14803 ( .A(M0_U3_U1_enc_tree_1__4__16_), .Y(n7348) );
  NAND2XL U14804 ( .A(n10731), .B(n10730), .Y(n7350) );
  OAI22XL U14805 ( .A0(n17092), .A1(n17086), .B0(n17099), .B1(n3022), .Y(
        n17095) );
  OAI2BB1XL U14806 ( .A0N(n16319), .A1N(n17087), .B0(n17073), .Y(n17094) );
  INVXL U14807 ( .A(M0_U4_U1_or2_tree_0__2__24_), .Y(M0_U4_U1_or2_inv_0__24_)
         );
  OR2XL U14808 ( .A(M0_U4_U1_or2_tree_0__2__16_), .B(
        M0_U4_U1_or2_tree_0__2__24_), .Y(n26149) );
  NOR2XL U14809 ( .A(n5397), .B(M0_a_12_), .Y(M0_U3_U1_enc_tree_0__1__18_) );
  INVXL U14810 ( .A(M0_U3_U1_or2_tree_0__2__24_), .Y(M0_U3_U1_or2_inv_0__24_)
         );
  OR2XL U14811 ( .A(M0_U3_U1_or2_tree_0__2__16_), .B(
        M0_U3_U1_or2_tree_0__2__24_), .Y(n26152) );
  INVXL U14812 ( .A(n12946), .Y(n12949) );
  INVXL U14813 ( .A(M3_U3_U1_enc_tree_1__4__16_), .Y(n12964) );
  AOI22XL U14814 ( .A0(n12948), .A1(n12947), .B0(n18804), .B1(n12949), .Y(
        n12953) );
  NAND2XL U14815 ( .A(n18800), .B(n12946), .Y(n12947) );
  OAI22XL U14816 ( .A0(n12965), .A1(n12942), .B0(n12941), .B1(
        M3_U3_U1_enc_tree_1__4__16_), .Y(n12963) );
  NOR2XL U14817 ( .A(n18822), .B(n12964), .Y(n12942) );
  INVXL U14818 ( .A(M3_U3_U1_enc_tree_2__4__16_), .Y(n12961) );
  OAI22X1 U14819 ( .A0(n17074), .A1(n16868), .B0(n16375), .B1(n16892), .Y(
        n16896) );
  OAI22X1 U14820 ( .A0(n16892), .A1(n17087), .B0(n16375), .B1(n5060), .Y(
        n16912) );
  CMPR32X1 U14821 ( .A(n16907), .B(n16906), .C(n16905), .CO(n16927), .S(n16901) );
  OAI22XL U14822 ( .A0(n16962), .A1(n3211), .B0(n16960), .B1(n16909), .Y(
        n16924) );
  OAI22XL U14823 ( .A0(n17060), .A1(n16904), .B0(n17061), .B1(n16923), .Y(
        n16919) );
  OAI21X1 U14824 ( .A0(n16319), .A1(n5067), .B0(n5065), .Y(n16920) );
  OAI21X1 U14825 ( .A0(n17044), .A1(n16375), .B0(n5063), .Y(n17043) );
  OAI22XL U14826 ( .A0(n17060), .A1(n17039), .B0(n17061), .B1(n17038), .Y(
        n17056) );
  XOR2XL U14827 ( .A(n22640), .B(n11209), .Y(M6_mult_x_15_n1142) );
  XOR2XL U14828 ( .A(n22792), .B(n3058), .Y(M6_mult_x_15_n1070) );
  XOR2XL U14829 ( .A(n22907), .B(n3053), .Y(M6_mult_x_15_n1166) );
  XOR2XL U14830 ( .A(n22756), .B(n3119), .Y(M6_mult_x_15_n1046) );
  OAI21XL U14831 ( .A0(n16734), .A1(n16735), .B0(n16733), .Y(n5735) );
  AOI22XL U14832 ( .A0(n21166), .A1(sigma12[0]), .B0(in_valid_t), .B1(w2[64]), 
        .Y(n15943) );
  NAND2X1 U14833 ( .A(in_valid_t), .B(w2[86]), .Y(n6018) );
  NAND2X1 U14834 ( .A(n21166), .B(sigma12[22]), .Y(n6019) );
  NAND2X1 U14835 ( .A(n5770), .B(data[118]), .Y(n6020) );
  INVXL U14836 ( .A(M5_U3_U1_enc_tree_3__3__16_), .Y(n17268) );
  INVXL U14837 ( .A(M5_U3_U1_enc_tree_1__4__16_), .Y(n17287) );
  AOI22XL U14838 ( .A0(n17271), .A1(n17270), .B0(n18804), .B1(n17272), .Y(
        n17276) );
  NAND2XL U14839 ( .A(n18800), .B(n17269), .Y(n17270) );
  INVXL U14840 ( .A(n17272), .Y(n17269) );
  INVXL U14841 ( .A(M5_U3_U1_enc_tree_2__4__16_), .Y(n17284) );
  NAND2X1 U14842 ( .A(in_valid_t), .B(w2[34]), .Y(n5050) );
  INVXL U14843 ( .A(M4_U4_U1_enc_tree_1__2__12_), .Y(
        M3_U4_U1_enc_tree_1__3__8_) );
  INVXL U14844 ( .A(M4_U3_U1_enc_tree_1__2__12_), .Y(
        M4_U3_U1_enc_tree_1__3__8_) );
  OR2XL U14845 ( .A(M4_U3_U1_or2_tree_1__2__16_), .B(
        M4_U3_U1_or2_tree_1__2__24_), .Y(n26150) );
  INVXL U14846 ( .A(n18822), .Y(n12941) );
  AOI21XL U14847 ( .A0(n22891), .A1(n3218), .B0(n22550), .Y(n22551) );
  OAI2BB1XL U14848 ( .A0N(n11071), .A1N(n22708), .B0(n22709), .Y(n22550) );
  INVXL U14849 ( .A(n22547), .Y(n22548) );
  NAND2XL U14850 ( .A(n10796), .B(n10795), .Y(n11221) );
  NAND2XL U14851 ( .A(w2[33]), .B(n23973), .Y(n10796) );
  NAND2XL U14852 ( .A(w2[65]), .B(valid[0]), .Y(n10795) );
  INVXL U14853 ( .A(n11222), .Y(n11207) );
  NAND2XL U14854 ( .A(n10753), .B(n10752), .Y(n11216) );
  NAND2XL U14855 ( .A(w2[37]), .B(n23973), .Y(n10753) );
  NAND2XL U14856 ( .A(w2[69]), .B(valid[0]), .Y(n10752) );
  NAND2XL U14857 ( .A(n10780), .B(n10779), .Y(n11219) );
  NAND2XL U14858 ( .A(w2[35]), .B(n23973), .Y(n10780) );
  NAND2XL U14859 ( .A(w2[67]), .B(valid[0]), .Y(n10779) );
  NAND2XL U14860 ( .A(w2[34]), .B(n23973), .Y(n10778) );
  NAND2XL U14861 ( .A(w2[66]), .B(valid[0]), .Y(n10777) );
  AOI2BB1XL U14862 ( .A0N(n11168), .A1N(n11167), .B0(n11166), .Y(n11449) );
  AOI2BB1XL U14863 ( .A0N(n11165), .A1N(n11164), .B0(n11163), .Y(n11167) );
  AOI2BB1XL U14864 ( .A0N(n11162), .A1N(n11161), .B0(n11160), .Y(n11164) );
  AOI2BB1XL U14865 ( .A0N(n11159), .A1N(n11158), .B0(n22867), .Y(n11161) );
  NOR2XL U14866 ( .A(n11067), .B(n22582), .Y(n11069) );
  NAND2XL U14867 ( .A(n22586), .B(n11065), .Y(n11067) );
  AOI21XL U14868 ( .A0(n22891), .A1(n11071), .B0(n22708), .Y(n22494) );
  INVXL U14869 ( .A(n23152), .Y(n23073) );
  NOR2XL U14870 ( .A(n22505), .B(n11079), .Y(n21068) );
  NOR2XL U14871 ( .A(n22515), .B(n11077), .Y(n11078) );
  INVXL U14872 ( .A(n22517), .Y(n11077) );
  INVXL U14873 ( .A(n22506), .Y(n22570) );
  NAND2XL U14874 ( .A(w2[84]), .B(valid[0]), .Y(n11083) );
  NAND2XL U14875 ( .A(w2[52]), .B(n3501), .Y(n11084) );
  OAI21XL U14876 ( .A0(n16149), .A1(n16148), .B0(n16147), .Y(n4832) );
  XNOR2XL U14877 ( .A(n3203), .B(M3_mult_x_15_b_20_), .Y(n16279) );
  INVX1 U14878 ( .A(n19374), .Y(n19820) );
  INVXL U14879 ( .A(n19557), .Y(n19598) );
  INVXL U14880 ( .A(n19563), .Y(n19736) );
  INVXL U14881 ( .A(n19538), .Y(n19551) );
  INVX1 U14882 ( .A(n19445), .Y(n19922) );
  INVXL U14883 ( .A(n20411), .Y(n20434) );
  NAND2XL U14884 ( .A(n3040), .B(n8357), .Y(n8358) );
  NOR2X2 U14885 ( .A(n7236), .B(n7257), .Y(n7320) );
  NAND2XL U14886 ( .A(n6953), .B(n6952), .Y(n5134) );
  NAND2XL U14887 ( .A(n19424), .B(n19914), .Y(n19916) );
  AOI21XL U14888 ( .A0(n19921), .A1(n19952), .B0(n3164), .Y(n19920) );
  OAI22XL U14889 ( .A0(n19928), .A1(n3100), .B0(n3041), .B1(n19927), .Y(n19943) );
  OAI22XL U14890 ( .A0(n7829), .A1(n7800), .B0(n7828), .B1(n25872), .Y(n7736)
         );
  OAI22XL U14891 ( .A0(n4642), .A1(n23219), .B0(n7712), .B1(n7711), .Y(n7737)
         );
  CMPR32X1 U14892 ( .A(n7691), .B(n7690), .C(n7689), .CO(n7709), .S(n7692) );
  INVXL U14893 ( .A(n25875), .Y(n7691) );
  OAI22XL U14894 ( .A0(n4642), .A1(n7647), .B0(n7696), .B1(n7712), .Y(n7690)
         );
  OAI22XL U14895 ( .A0(n7829), .A1(n25873), .B0(n7828), .B1(n7800), .Y(n7715)
         );
  NAND2XL U14896 ( .A(n5124), .B(n7695), .Y(n5110) );
  NAND2X1 U14897 ( .A(n9368), .B(n9367), .Y(n5390) );
  OAI22XL U14898 ( .A0(n10517), .A1(n10495), .B0(n10533), .B1(n10494), .Y(
        n10510) );
  INVXL U14899 ( .A(n10515), .Y(n10516) );
  OAI22XL U14900 ( .A0(n10660), .A1(M2_mult_x_15_n1669), .B0(n10659), .B1(
        M2_mult_x_15_n1668), .Y(n10550) );
  NOR2X1 U14901 ( .A(n5257), .B(n10554), .Y(n5256) );
  AND2XL U14902 ( .A(n10250), .B(M2_U4_U1_enc_tree_3__3__24_), .Y(n10256) );
  INVXL U14903 ( .A(M2_U4_U1_enc_tree_3__3__16_), .Y(n10250) );
  NAND2XL U14904 ( .A(n10249), .B(M2_U3_U1_enc_tree_3__3__24_), .Y(n10252) );
  INVXL U14905 ( .A(M2_U3_U1_enc_tree_3__3__16_), .Y(n10249) );
  INVXL U14906 ( .A(n10252), .Y(n10257) );
  INVXL U14907 ( .A(M2_U4_U1_enc_tree_1__2__12_), .Y(
        M2_U4_U1_enc_tree_1__3__8_) );
  OR2XL U14908 ( .A(M2_U4_U1_or2_tree_1__2__16_), .B(
        M2_U4_U1_or2_tree_1__2__24_), .Y(n26153) );
  OR2XL U14909 ( .A(M2_U3_U1_or2_tree_1__2__16_), .B(
        M2_U3_U1_or2_tree_1__2__24_), .Y(n26205) );
  INVXL U14910 ( .A(M2_U4_U1_enc_tree_2__4__16_), .Y(n10266) );
  INVXL U14911 ( .A(M2_U3_U1_enc_tree_2__4__16_), .Y(n10267) );
  INVXL U14912 ( .A(M2_U4_U1_enc_tree_1__4__16_), .Y(n10270) );
  INVXL U14913 ( .A(M2_U3_U1_enc_tree_1__4__16_), .Y(n10271) );
  INVXL U14914 ( .A(M2_U3_U1_enc_tree_0__4__16_), .Y(n10705) );
  OR2XL U14915 ( .A(M2_U3_U1_or2_tree_0__2__16_), .B(
        M2_U3_U1_or2_tree_0__2__24_), .Y(n26207) );
  INVXL U14916 ( .A(M2_U4_U1_enc_tree_0__4__16_), .Y(n10704) );
  INVXL U14917 ( .A(M2_U4_U1_enc_tree_0__2__12_), .Y(
        M2_U4_U1_enc_tree_0__3__8_) );
  OR2XL U14918 ( .A(M2_U4_U1_or2_tree_0__2__16_), .B(
        M2_U4_U1_or2_tree_0__2__24_), .Y(n26156) );
  NOR2X1 U14919 ( .A(n4890), .B(n12633), .Y(n4889) );
  OAI22X1 U14920 ( .A0(n12340), .A1(n11727), .B0(n12338), .B1(n2980), .Y(
        n11730) );
  OAI22XL U14921 ( .A0(n12352), .A1(n11830), .B0(n12222), .B1(n11746), .Y(
        n11810) );
  OAI22X1 U14922 ( .A0(n12759), .A1(n11813), .B0(n12760), .B1(n11812), .Y(
        n11856) );
  OAI22XL U14923 ( .A0(n12578), .A1(n12516), .B0(n12718), .B1(n12539), .Y(
        n12543) );
  OAI22X1 U14924 ( .A0(n12618), .A1(n12515), .B0(n12616), .B1(n5956), .Y(
        n12544) );
  OAI22XL U14925 ( .A0(n12717), .A1(n12539), .B0(n12718), .B1(n12555), .Y(
        n12558) );
  OAI22XL U14926 ( .A0(n12717), .A1(n12716), .B0(n12718), .B1(n12696), .Y(
        n12711) );
  CMPR32X1 U14927 ( .A(n18471), .B(n18470), .C(n18469), .CO(n18475), .S(n18454) );
  OAI22XL U14928 ( .A0(n18522), .A1(n18452), .B0(n3195), .B1(n18468), .Y(
        n18470) );
  CMPR32X1 U14929 ( .A(n12542), .B(n18447), .C(n18446), .CO(n18456), .S(n18441) );
  OAI22XL U14930 ( .A0(n18721), .A1(M3_mult_x_15_b_13_), .B0(n17512), .B1(
        n18611), .Y(n18447) );
  OAI22XL U14931 ( .A0(n12759), .A1(n12745), .B0(n12760), .B1(n12758), .Y(
        n12754) );
  CMPR32X1 U14932 ( .A(n18548), .B(n18547), .C(n18546), .CO(n18565), .S(n18557) );
  OAI22XL U14933 ( .A0(n18652), .A1(n18545), .B0(n18653), .B1(n18544), .Y(
        n18546) );
  OAI22XL U14934 ( .A0(n18659), .A1(n18543), .B0(n17832), .B1(n18542), .Y(
        n18547) );
  XOR2X1 U14935 ( .A(n18350), .B(n5878), .Y(n18377) );
  XOR2X1 U14936 ( .A(n18352), .B(n18351), .Y(n5878) );
  OAI22X1 U14937 ( .A0(n18111), .A1(n17695), .B0(n18504), .B1(n17602), .Y(
        n17677) );
  OAI21XL U14938 ( .A0(n13442), .A1(n13441), .B0(n13440), .Y(n5260) );
  CMPR32X1 U14939 ( .A(n13680), .B(n13679), .C(n13678), .CO(n13750), .S(n13746) );
  OAI22XL U14940 ( .A0(n13653), .A1(n14198), .B0(n13618), .B1(n14208), .Y(
        n13678) );
  OAI22XL U14941 ( .A0(n13649), .A1(n14227), .B0(n13616), .B1(n14249), .Y(
        n13680) );
  OAI22XL U14942 ( .A0(n13654), .A1(n13972), .B0(n13617), .B1(n13971), .Y(
        n13679) );
  CMPR32X1 U14943 ( .A(n13660), .B(n13659), .C(n13658), .CO(n13707), .S(n13745) );
  OAI22XL U14944 ( .A0(n13666), .A1(n14120), .B0(n13619), .B1(n14121), .Y(
        n13660) );
  NAND2BXL U14945 ( .AN(n13049), .B(n23173), .Y(n13511) );
  INVXL U14946 ( .A(M1_U4_U1_enc_tree_3__3__16_), .Y(n14366) );
  INVXL U14947 ( .A(n14368), .Y(n14372) );
  INVXL U14948 ( .A(M1_U3_U1_enc_tree_1__4__16_), .Y(n14386) );
  INVXL U14949 ( .A(M1_U4_U1_enc_tree_1__4__16_), .Y(n14385) );
  AOI22XL U14950 ( .A0(n14370), .A1(n14369), .B0(n14371), .B1(n14372), .Y(
        n14376) );
  NAND2XL U14951 ( .A(n14368), .B(n14367), .Y(n14369) );
  INVXL U14952 ( .A(n14371), .Y(n14367) );
  NOR2XL U14953 ( .A(n14379), .B(n14378), .Y(n14377) );
  OAI22XL U14954 ( .A0(n14363), .A1(n14387), .B0(M1_U3_U1_enc_tree_1__4__16_), 
        .B1(M1_U4_U1_enc_tree_1__4__16_), .Y(n14392) );
  NOR2XL U14955 ( .A(n14386), .B(n14385), .Y(n14363) );
  INVXL U14956 ( .A(M1_U4_U1_enc_tree_2__4__16_), .Y(n14389) );
  INVXL U14957 ( .A(M1_U3_U1_enc_tree_2__4__16_), .Y(n14390) );
  INVXL U14958 ( .A(M1_U4_U1_enc_tree_0__4__16_), .Y(n14478) );
  INVXL U14959 ( .A(M1_U4_U1_enc_tree_0__2__12_), .Y(
        M1_U4_U1_enc_tree_0__3__8_) );
  INVXL U14960 ( .A(M1_U3_U1_enc_tree_0__4__16_), .Y(n14479) );
  OR2XL U14961 ( .A(M1_U3_U1_or2_tree_0__2__16_), .B(
        M1_U3_U1_or2_tree_0__2__24_), .Y(n26209) );
  OAI22X1 U14962 ( .A0(n18624), .A1(n17747), .B0(n18625), .B1(n17779), .Y(
        n17789) );
  CMPR32X1 U14963 ( .A(n18519), .B(n18518), .C(n18517), .CO(n18562), .S(n18584) );
  OAI22XL U14964 ( .A0(n18652), .A1(n17834), .B0(n18653), .B1(n18545), .Y(
        n18517) );
  OAI22XL U14965 ( .A0(n18659), .A1(n17833), .B0(n17832), .B1(n18543), .Y(
        n18518) );
  ADDFX2 U14966 ( .A(n14207), .B(n14206), .CI(n14205), .CO(n14223), .S(n14218)
         );
  OAI22XL U14967 ( .A0(n14148), .A1(n14208), .B0(n14198), .B1(M1_b_15_), .Y(
        n14193) );
  OAI22XL U14968 ( .A0(n14115), .A1(n14249), .B0(n14159), .B1(n14250), .Y(
        n14147) );
  CMPR32X1 U14969 ( .A(n12642), .B(n12641), .C(n12640), .CO(n12659), .S(n12651) );
  OAI22XL U14970 ( .A0(n12715), .A1(n12639), .B0(n12746), .B1(n12638), .Y(
        n12640) );
  OAI22X1 U14971 ( .A0(n12746), .A1(n11985), .B0(n12715), .B1(n4906), .Y(
        n11977) );
  NOR2X2 U14972 ( .A(n3415), .B(n12820), .Y(n6111) );
  INVXL U14973 ( .A(n12815), .Y(n12816) );
  OAI21XL U14974 ( .A0(n5461), .A1(n18213), .B0(n18212), .Y(n18214) );
  NAND2XL U14975 ( .A(n18267), .B(n18261), .Y(n18269) );
  OAI22XL U14976 ( .A0(n18624), .A1(n18604), .B0(n18625), .B1(n18603), .Y(
        n18621) );
  CMPR32X1 U14977 ( .A(n3107), .B(n18486), .C(n18485), .CO(n18600), .S(n18476)
         );
  OAI22XL U14978 ( .A0(n18721), .A1(n3198), .B0(n17512), .B1(n3021), .Y(n18486) );
  OAI22XL U14979 ( .A0(n18522), .A1(n18468), .B0(n3195), .B1(n18467), .Y(
        n18485) );
  OAI2BB1XL U14980 ( .A0N(n3195), .A1N(n18483), .B0(n18468), .Y(n18605) );
  CMPR32X1 U14981 ( .A(n18480), .B(n18479), .C(n18478), .CO(n18614), .S(n18489) );
  OAI22XL U14982 ( .A0(n18624), .A1(n18462), .B0(n18625), .B1(n18484), .Y(
        n18478) );
  OAI22XL U14983 ( .A0(n18652), .A1(n18461), .B0(n18653), .B1(n18481), .Y(
        n18479) );
  OAI22XL U14984 ( .A0(n14233), .A1(n14282), .B0(n14252), .B1(n14251), .Y(
        n14244) );
  OAI22XL U14985 ( .A0(n14232), .A1(n6191), .B0(n14253), .B1(n14298), .Y(
        n14245) );
  ADDFX2 U14986 ( .A(n14226), .B(n14225), .CI(n14224), .CO(n14242), .S(n14237)
         );
  OAI22XL U14987 ( .A0(n14214), .A1(n14249), .B0(n14250), .B1(n14228), .Y(
        n14226) );
  NAND2XL U14988 ( .A(n13787), .B(n13786), .Y(n13788) );
  INVXL U14989 ( .A(n14307), .Y(n14301) );
  OAI22XL U14990 ( .A0(n6191), .A1(n23173), .B0(n14298), .B1(n14290), .Y(
        n14299) );
  OAI22XL U14991 ( .A0(n2993), .A1(n14306), .B0(n14289), .B1(n14357), .Y(
        n14300) );
  AOI2BB2XL U14992 ( .B0(n19724), .B1(n19542), .A0N(n19693), .A1N(n19542), .Y(
        n19694) );
  INVXL U14993 ( .A(n8742), .Y(n8743) );
  INVXL U14994 ( .A(n8745), .Y(n8733) );
  NAND2XL U14995 ( .A(n8741), .B(n8746), .Y(n8735) );
  NAND2XL U14996 ( .A(n8700), .B(n8699), .Y(n8737) );
  AOI21XL U14997 ( .A0(n8860), .A1(n8729), .B0(n8720), .Y(n8721) );
  INVXL U14998 ( .A(n8728), .Y(n8720) );
  NAND2XL U14999 ( .A(n8853), .B(n8729), .Y(n8722) );
  NAND2XL U15000 ( .A(n8853), .B(n8851), .Y(n8708) );
  INVXL U15001 ( .A(n8774), .Y(n8853) );
  AOI21XL U15002 ( .A0(n8771), .A1(n8823), .B0(n3155), .Y(n8770) );
  AOI21XL U15003 ( .A0(n8792), .A1(n8823), .B0(n3155), .Y(n8791) );
  AOI21XL U15004 ( .A0(n8787), .A1(n8823), .B0(n3155), .Y(n8786) );
  AOI21XL U15005 ( .A0(n8802), .A1(n8823), .B0(n3155), .Y(n8801) );
  OAI22XL U15006 ( .A0(n8804), .A1(n3017), .B0(n3040), .B1(n8803), .Y(n8816)
         );
  OAI22XL U15007 ( .A0(n8607), .A1(n4591), .B0(n8606), .B1(n8605), .Y(n8609)
         );
  OAI22XL U15008 ( .A0(n8451), .A1(n3087), .B0(n3157), .B1(n8448), .Y(n8613)
         );
  NAND2XL U15009 ( .A(n8696), .B(n8695), .Y(n8750) );
  INVXL U15010 ( .A(n8719), .Y(n8729) );
  NOR2XL U15011 ( .A(n9017), .B(n20390), .Y(n9018) );
  INVXL U15012 ( .A(n20199), .Y(n20175) );
  INVXL U15013 ( .A(n20046), .Y(n19889) );
  NOR2XL U15014 ( .A(n19888), .B(n20048), .Y(n19891) );
  INVXL U15015 ( .A(n20047), .Y(n19888) );
  NAND2XL U15016 ( .A(n19767), .B(n19766), .Y(n20054) );
  INVXL U15017 ( .A(n20053), .Y(n20044) );
  NAND2XL U15018 ( .A(n20023), .B(n20022), .Y(n20024) );
  INVXL U15019 ( .A(n20021), .Y(n20023) );
  INVXL U15020 ( .A(n15667), .Y(n15509) );
  NOR2XL U15021 ( .A(n15508), .B(n15669), .Y(n15511) );
  INVXL U15022 ( .A(n15668), .Y(n15508) );
  INVXL U15023 ( .A(n15491), .Y(n15492) );
  OAI22XL U15024 ( .A0(n21776), .A1(n3042), .B0(n23116), .B1(n21195), .Y(
        n21811) );
  INVXL U15025 ( .A(n21626), .Y(n21810) );
  NAND2XL U15026 ( .A(n21178), .B(n21177), .Y(n21625) );
  NAND3XL U15027 ( .A(cs[0]), .B(cs[1]), .C(target_temp[3]), .Y(n21177) );
  NAND2XL U15028 ( .A(n21628), .B(n21977), .Y(n21518) );
  NAND2XL U15029 ( .A(n21628), .B(n21997), .Y(n21512) );
  NAND2XL U15030 ( .A(n21628), .B(n21992), .Y(n21510) );
  NAND2XL U15031 ( .A(n21560), .B(n3095), .Y(n21712) );
  NAND2XL U15032 ( .A(n21331), .B(w1[13]), .Y(n21252) );
  INVXL U15033 ( .A(n21457), .Y(n21871) );
  NAND2XL U15034 ( .A(n21331), .B(w1[11]), .Y(n21237) );
  INVXL U15035 ( .A(n21475), .Y(n21853) );
  INVXL U15036 ( .A(n21604), .Y(n21617) );
  INVXL U15037 ( .A(n21460), .Y(n21876) );
  NAND2XL U15038 ( .A(n21244), .B(n21243), .Y(n21552) );
  NAND3XL U15039 ( .A(cs[0]), .B(cs[1]), .C(y20[9]), .Y(n21243) );
  INVXL U15040 ( .A(n21470), .Y(n21553) );
  AOI2BB2XL U15041 ( .B0(n23116), .B1(n21656), .A0N(n23116), .A1N(n21657), .Y(
        n21701) );
  AOI2BB2XL U15042 ( .B0(n23116), .B1(n21639), .A0N(n21628), .A1N(n21640), .Y(
        n21700) );
  INVXL U15043 ( .A(n21513), .Y(n21902) );
  INVXL U15044 ( .A(n21456), .Y(n21863) );
  INVXL U15045 ( .A(n21554), .Y(n21579) );
  NAND2XL U15046 ( .A(n21186), .B(n21185), .Y(n21775) );
  INVXL U15047 ( .A(n21623), .Y(n21776) );
  AOI2BB2XL U15048 ( .B0(n23116), .B1(n21987), .A0N(n21628), .A1N(n21988), .Y(
        n21676) );
  INVXL U15049 ( .A(n21473), .Y(n21845) );
  INVXL U15050 ( .A(n21469), .Y(n21531) );
  INVXL U15051 ( .A(n21556), .Y(n21601) );
  NOR2XL U15052 ( .A(n21478), .B(n21481), .Y(n21484) );
  OAI21XL U15053 ( .A0(n21481), .A1(n21480), .B0(n21479), .Y(n21482) );
  NAND2XL U15054 ( .A(n21201), .B(n21626), .Y(n21202) );
  NAND2XL U15055 ( .A(n21200), .B(n21625), .Y(n21203) );
  NAND2XL U15056 ( .A(n21184), .B(n21189), .Y(n21199) );
  AOI21XL U15057 ( .A0(n21189), .A1(n6185), .B0(n21196), .Y(n21197) );
  AND2XL U15058 ( .A(n21194), .B(n21620), .Y(n6185) );
  NOR2XL U15059 ( .A(n21200), .B(n21625), .Y(n21179) );
  NAND2XL U15060 ( .A(n21220), .B(n21554), .Y(n21221) );
  NAND2XL U15061 ( .A(n21224), .B(n21556), .Y(n21227) );
  NAND2XL U15062 ( .A(n21266), .B(n21456), .Y(n21267) );
  NAND2XL U15063 ( .A(n21470), .B(n21260), .Y(n21263) );
  NAND2XL U15064 ( .A(n21274), .B(n21460), .Y(n21275) );
  NAND2XL U15065 ( .A(n21278), .B(n21461), .Y(n21281) );
  INVXL U15066 ( .A(n21552), .Y(n21260) );
  NAND2XL U15067 ( .A(n15645), .B(n15644), .Y(n15646) );
  INVXL U15068 ( .A(n15643), .Y(n15645) );
  INVXL U15069 ( .A(n15494), .Y(n15482) );
  NAND2XL U15070 ( .A(n15490), .B(n15495), .Y(n15484) );
  NAND2XL U15071 ( .A(n15449), .B(n15448), .Y(n15486) );
  AOI21XL U15072 ( .A0(n15610), .A1(n15609), .B0(n15608), .Y(n15611) );
  INVXL U15073 ( .A(n15604), .Y(n15607) );
  NAND2XL U15074 ( .A(n15603), .B(n15609), .Y(n15612) );
  NAND2XL U15075 ( .A(n15453), .B(n15452), .Y(n15477) );
  INVXL U15076 ( .A(n15468), .Y(n15478) );
  NAND2XL U15077 ( .A(n15046), .B(n15437), .Y(n15439) );
  OAI22XL U15078 ( .A0(n15441), .A1(n3101), .B0(n15008), .B1(n15440), .Y(
        n15454) );
  INVXL U15079 ( .A(n15530), .Y(n15610) );
  INVXL U15080 ( .A(n15523), .Y(n15603) );
  NAND2XL U15081 ( .A(n15046), .B(n15458), .Y(n15460) );
  OAI22XL U15082 ( .A0(n15462), .A1(n3101), .B0(n15008), .B1(n15461), .Y(
        n15463) );
  NAND2XL U15083 ( .A(n21792), .B(n22086), .Y(n22087) );
  NAND2XL U15084 ( .A(n22082), .B(n22081), .Y(n22083) );
  INVXL U15085 ( .A(n22080), .Y(n22082) );
  INVXL U15086 ( .A(n22104), .Y(n21949) );
  NOR2XL U15087 ( .A(n21948), .B(n22106), .Y(n21951) );
  INVXL U15088 ( .A(n22105), .Y(n21948) );
  NAND2XL U15089 ( .A(n21834), .B(n21833), .Y(n21953) );
  NAND2XL U15090 ( .A(n21893), .B(n21892), .Y(n21917) );
  INVXL U15091 ( .A(n21908), .Y(n21918) );
  OAI21XL U15092 ( .A0(n21854), .A1(n21981), .B0(n21980), .Y(n22002) );
  AOI21XL U15093 ( .A0(n21981), .A1(n3222), .B0(n21849), .Y(n21980) );
  OAI22XL U15094 ( .A0(n21983), .A1(n21429), .B0(n3020), .B1(n21342), .Y(
        n22001) );
  AOI21XL U15095 ( .A0(n21986), .A1(n3222), .B0(n21849), .Y(n21985) );
  NAND2XL U15096 ( .A(n21506), .B(n21984), .Y(n21986) );
  OAI22XL U15097 ( .A0(n21988), .A1(n3042), .B0(n3020), .B1(n21343), .Y(n22003) );
  AOI21XL U15098 ( .A0(n21976), .A1(n3222), .B0(n21849), .Y(n21975) );
  OAI22XL U15099 ( .A0(n21978), .A1(n21429), .B0(n3020), .B1(n21338), .Y(
        n21999) );
  OAI21XL U15100 ( .A0(n21854), .A1(n21960), .B0(n21959), .Y(n21965) );
  AOI21XL U15101 ( .A0(n21960), .A1(n3222), .B0(n21849), .Y(n21959) );
  NAND2XL U15102 ( .A(n21506), .B(n21958), .Y(n21960) );
  OAI22XL U15103 ( .A0(n21962), .A1(n21429), .B0(n3020), .B1(n21337), .Y(
        n21964) );
  AOI21XL U15104 ( .A0(n21991), .A1(n3222), .B0(n21849), .Y(n21990) );
  OAI22XL U15105 ( .A0(n21993), .A1(n3042), .B0(n3020), .B1(n21350), .Y(n22005) );
  INVXL U15106 ( .A(n21934), .Y(n21922) );
  NAND2XL U15107 ( .A(n21930), .B(n21935), .Y(n21924) );
  NAND2XL U15108 ( .A(n21889), .B(n21888), .Y(n21926) );
  AOI21XL U15109 ( .A0(n22048), .A1(n21918), .B0(n21909), .Y(n21910) );
  INVXL U15110 ( .A(n21917), .Y(n21909) );
  NAND2XL U15111 ( .A(n22041), .B(n21918), .Y(n21911) );
  NAND2XL U15112 ( .A(n21895), .B(n21894), .Y(n21913) );
  NAND2XL U15113 ( .A(n22041), .B(n22039), .Y(n21897) );
  NAND2XL U15114 ( .A(n21904), .B(n21903), .Y(n22043) );
  NAND4XL U15115 ( .A(n22301), .B(n22203), .C(n22202), .D(n22305), .Y(n22204)
         );
  NAND2XL U15116 ( .A(n21887), .B(n21886), .Y(n21934) );
  INVXL U15117 ( .A(n21921), .Y(n21935) );
  OAI21XL U15118 ( .A0(n21938), .A1(n21944), .B0(n21939), .Y(n21931) );
  INVXL U15119 ( .A(n21930), .Y(n21933) );
  AOI211XL U15120 ( .A0(n8972), .A1(n8971), .B0(n20453), .C0(n20454), .Y(n8974) );
  AOI211XL U15121 ( .A0(n8967), .A1(n8966), .B0(n20435), .C0(n20436), .Y(n8970) );
  OAI21XL U15122 ( .A0(n17065), .A1(n17067), .B0(n17066), .Y(n5094) );
  NOR2XL U15123 ( .A(M6_mult_x_15_n509), .B(M6_mult_x_15_n517), .Y(n10990) );
  XNOR2X1 U15124 ( .A(n11694), .B(n11693), .Y(n4956) );
  NAND2XL U15125 ( .A(n11351), .B(n11000), .Y(n11006) );
  XOR2XL U15126 ( .A(n22536), .B(n3119), .Y(M6_mult_x_15_n1034) );
  INVXL U15127 ( .A(n23102), .Y(M6_mult_x_15_n1010) );
  XOR2XL U15128 ( .A(n22525), .B(n3119), .Y(M6_mult_x_15_n1033) );
  XOR2XL U15129 ( .A(n22538), .B(n3119), .Y(M6_mult_x_15_n1032) );
  XOR2XL U15130 ( .A(n22615), .B(n11209), .Y(M6_mult_x_15_n1140) );
  XOR2XL U15131 ( .A(n22617), .B(n3055), .Y(M6_mult_x_15_n1115) );
  NAND2XL U15132 ( .A(M6_mult_x_15_n528), .B(M6_mult_x_15_n537), .Y(n11345) );
  NOR2XL U15133 ( .A(n11124), .B(n11126), .Y(n11108) );
  XOR2XL U15134 ( .A(n22545), .B(n3058), .Y(M6_mult_x_15_n1061) );
  XOR2XL U15135 ( .A(n22510), .B(n3058), .Y(M6_mult_x_15_n1060) );
  INVXL U15136 ( .A(n10997), .Y(n11351) );
  NOR2BXL U15137 ( .AN(n11207), .B(n10798), .Y(n22897) );
  AOI222XL U15138 ( .A0(n22953), .A1(n3218), .B0(n22897), .B1(n23089), .C0(
        n22952), .C1(n11074), .Y(n22623) );
  XOR2XL U15139 ( .A(n22742), .B(n3058), .Y(M6_mult_x_15_n1074) );
  XOR2XL U15140 ( .A(n22678), .B(n3056), .Y(M6_mult_x_15_n1098) );
  XOR2XL U15141 ( .A(n22858), .B(n3119), .Y(M6_mult_x_15_n1050) );
  XOR2XL U15142 ( .A(n22692), .B(n3056), .Y(M6_mult_x_15_n1097) );
  XOR2XL U15143 ( .A(n22733), .B(n3119), .Y(M6_mult_x_15_n1049) );
  XOR2XL U15144 ( .A(n22817), .B(n3058), .Y(M6_mult_x_15_n1073) );
  XOR2XL U15145 ( .A(n22819), .B(n3054), .Y(M6_mult_x_15_n1145) );
  XOR2XL U15146 ( .A(n22811), .B(n3053), .Y(M6_mult_x_15_n1169) );
  XOR2XL U15147 ( .A(n11257), .B(n11256), .Y(n11258) );
  NAND2XL U15148 ( .A(n11258), .B(n11265), .Y(n11260) );
  AOI211XL U15149 ( .A0(n11139), .A1(n11138), .B0(n11166), .C0(n11168), .Y(
        n11270) );
  NOR2BXL U15150 ( .AN(n11252), .B(n11251), .Y(n11265) );
  XOR2XL U15151 ( .A(n7335), .B(n7334), .Y(n7336) );
  INVXL U15152 ( .A(n7339), .Y(n7344) );
  INVXL U15153 ( .A(n7340), .Y(n7343) );
  OAI22XL U15154 ( .A0(n7350), .A1(n7327), .B0(M0_U4_U1_enc_tree_1__4__16_), 
        .B1(M0_U3_U1_enc_tree_1__4__16_), .Y(n7355) );
  NOR2XL U15155 ( .A(n7349), .B(n7348), .Y(n7327) );
  XOR2XL U15156 ( .A(n7353), .B(n7352), .Y(n7354) );
  NAND2XL U15157 ( .A(n7339), .B(n7340), .Y(n7347) );
  XOR2XL U15158 ( .A(n7351), .B(n7350), .Y(n7357) );
  XOR2XL U15159 ( .A(n7349), .B(n7348), .Y(n7351) );
  AND2X1 U15160 ( .A(n6719), .B(n6718), .Y(n6720) );
  NAND2X1 U15161 ( .A(n6712), .B(n6713), .Y(n5623) );
  OAI21X1 U15162 ( .A0(n5550), .A1(n6675), .B0(n6674), .Y(n5549) );
  NOR2X1 U15163 ( .A(n5552), .B(n6675), .Y(n5551) );
  OAI22XL U15164 ( .A0(n17092), .A1(n3022), .B0(n17099), .B1(n6014), .Y(n17100) );
  OAI22XL U15165 ( .A0(n17148), .A1(M3_mult_x_15_b_21_), .B0(n17147), .B1(
        n3202), .Y(n17101) );
  NOR2XL U15166 ( .A(n18810), .B(n12955), .Y(n12954) );
  XOR2XL U15167 ( .A(n12951), .B(n12950), .Y(n12952) );
  XNOR2XL U15168 ( .A(n18804), .B(n12949), .Y(n12950) );
  INVXL U15169 ( .A(n12948), .Y(n12951) );
  INVXL U15170 ( .A(n12953), .Y(n12957) );
  XNOR2XL U15171 ( .A(n18822), .B(n12964), .Y(n12966) );
  NAND2XL U15172 ( .A(n12953), .B(n12954), .Y(n12960) );
  XOR2XL U15173 ( .A(n12963), .B(n12962), .Y(n12968) );
  XOR2XL U15174 ( .A(n18818), .B(n12961), .Y(n12962) );
  INVXL U15175 ( .A(M3_U3_U1_enc_tree_0__4__16_), .Y(n13031) );
  INVXL U15176 ( .A(M3_U3_U1_enc_tree_0__2__12_), .Y(
        M3_U3_U1_enc_tree_0__3__8_) );
  OR2XL U15177 ( .A(M3_U3_U1_or2_tree_0__2__16_), .B(
        M3_U3_U1_or2_tree_0__2__24_), .Y(n26158) );
  XOR2XL U15178 ( .A(n22626), .B(n3053), .Y(M6_mult_x_15_n1167) );
  OAI22XL U15179 ( .A0(n18652), .A1(n18623), .B0(n18653), .B1(n18638), .Y(
        n18633) );
  OAI22XL U15180 ( .A0(n18659), .A1(n18635), .B0(n17832), .B1(n18651), .Y(
        n18650) );
  OAI22XL U15181 ( .A0(n18659), .A1(n18651), .B0(n17832), .B1(n25883), .Y(
        n18662) );
  INVXL U15182 ( .A(n18967), .Y(n18701) );
  NOR2XL U15183 ( .A(n18810), .B(n17278), .Y(n17277) );
  XOR2XL U15184 ( .A(n17274), .B(n17273), .Y(n17275) );
  XNOR2XL U15185 ( .A(n18804), .B(n17272), .Y(n17273) );
  INVXL U15186 ( .A(n17271), .Y(n17274) );
  INVXL U15187 ( .A(n17276), .Y(n17280) );
  XNOR2XL U15188 ( .A(n18822), .B(n17287), .Y(n17289) );
  NAND2XL U15189 ( .A(n17276), .B(n17277), .Y(n17283) );
  XOR2XL U15190 ( .A(n17286), .B(n17285), .Y(n17291) );
  XOR2XL U15191 ( .A(n18818), .B(n17284), .Y(n17285) );
  AOI22XL U15192 ( .A0(n5480), .A1(sigma11[0]), .B0(in_valid_t), .B1(w2[32]), 
        .Y(n17479) );
  INVXL U15193 ( .A(M3_mult_x_15_b_17_), .Y(M4_U4_U1_or2_inv_0__14_) );
  INVXL U15194 ( .A(M3_mult_x_15_b_21_), .Y(M4_U4_U1_or2_inv_0__10_) );
  INVXL U15195 ( .A(M4_U3_U1_enc_tree_1__4__16_), .Y(n18821) );
  AOI22XL U15196 ( .A0(n18802), .A1(n18801), .B0(n18804), .B1(n18803), .Y(
        n18808) );
  NAND2XL U15197 ( .A(n18800), .B(n18799), .Y(n18801) );
  INVXL U15198 ( .A(n18803), .Y(n18799) );
  OAI22XL U15199 ( .A0(n18823), .A1(n18795), .B0(n12941), .B1(
        M4_U3_U1_enc_tree_1__4__16_), .Y(n18820) );
  NOR2XL U15200 ( .A(n18822), .B(n18821), .Y(n18795) );
  INVXL U15201 ( .A(M4_U3_U1_enc_tree_2__4__16_), .Y(n18817) );
  NAND2XL U15202 ( .A(n10969), .B(n10965), .Y(n11004) );
  INVXL U15203 ( .A(n23099), .Y(M6_mult_x_15_n1008) );
  XOR2XL U15204 ( .A(n22552), .B(n3119), .Y(M6_mult_x_15_n1031) );
  NOR2BXL U15205 ( .AN(n11449), .B(n11453), .Y(n11450) );
  INVXL U15206 ( .A(n22891), .Y(n22522) );
  XOR2XL U15207 ( .A(n22495), .B(n3119), .Y(M6_mult_x_15_n1030) );
  INVXL U15208 ( .A(n23092), .Y(M6_mult_x_15_n1007) );
  OAI2BB1XL U15209 ( .A0N(n11071), .A1N(n23093), .B0(n23073), .Y(n23074) );
  INVXL U15210 ( .A(n10964), .Y(n10953) );
  INVXL U15211 ( .A(n10968), .Y(n10954) );
  AOI21XL U15212 ( .A0(n11012), .A1(n11011), .B0(n11010), .Y(n11013) );
  INVXL U15213 ( .A(n11009), .Y(n11010) );
  INVXL U15214 ( .A(n11008), .Y(n11012) );
  NAND2XL U15215 ( .A(n11003), .B(n11011), .Y(n11014) );
  NOR2XL U15216 ( .A(n11004), .B(n11014), .Y(n11017) );
  NAND2XL U15217 ( .A(n11005), .B(n11017), .Y(n11020) );
  NOR2XL U15218 ( .A(n11036), .B(n11357), .Y(n11007) );
  AOI21XL U15219 ( .A0(n10942), .A1(n11039), .B0(n10941), .Y(n10984) );
  AOI21XL U15220 ( .A0(n10987), .A1(n10944), .B0(n10943), .Y(n10945) );
  NAND2XL U15221 ( .A(n10942), .B(n11038), .Y(n10985) );
  NAND2XL U15222 ( .A(n19455), .B(n19383), .Y(n19174) );
  INVXL U15223 ( .A(n19384), .Y(n19455) );
  INVXL U15224 ( .A(n9028), .Y(n9002) );
  INVXL U15225 ( .A(n20436), .Y(n20389) );
  NAND2XL U15226 ( .A(n3067), .B(n20439), .Y(n20388) );
  INVXL U15227 ( .A(n20432), .Y(n20387) );
  NAND2XL U15228 ( .A(n3067), .B(n20435), .Y(n20386) );
  NOR2XL U15229 ( .A(n3124), .B(n20445), .Y(n20446) );
  INVXL U15230 ( .A(n20443), .Y(n20444) );
  INVXL U15231 ( .A(n20435), .Y(n20438) );
  NAND2XL U15232 ( .A(n3067), .B(n20436), .Y(n20437) );
  INVXL U15233 ( .A(n20449), .Y(n20452) );
  INVXL U15234 ( .A(n9006), .Y(n9011) );
  INVXL U15235 ( .A(n20008), .Y(n19966) );
  INVXL U15236 ( .A(n10430), .Y(n5183) );
  NOR2X1 U15237 ( .A(n10228), .B(n10195), .Y(n10234) );
  AOI21XL U15238 ( .A0(n10233), .A1(n10192), .B0(n10191), .Y(n10193) );
  INVXL U15239 ( .A(n15629), .Y(n15587) );
  INVXL U15240 ( .A(n15580), .Y(n15622) );
  NAND3XL U15241 ( .A(n15861), .B(n15872), .C(n24871), .Y(n15771) );
  INVXL U15242 ( .A(n10648), .Y(n10649) );
  AND2X2 U15243 ( .A(n10052), .B(n10051), .Y(n5138) );
  NOR2XL U15244 ( .A(n10032), .B(n10039), .Y(n10040) );
  OAI22X1 U15245 ( .A0(n10046), .A1(n10045), .B0(n5179), .B1(n5178), .Y(n10050) );
  INVXL U15246 ( .A(n10255), .Y(n10259) );
  XNOR2XL U15247 ( .A(n10257), .B(n10256), .Y(n10258) );
  AOI22XL U15248 ( .A0(n10255), .A1(n10253), .B0(n10256), .B1(n10257), .Y(
        n10263) );
  NAND2XL U15249 ( .A(n10252), .B(n10251), .Y(n10253) );
  INVXL U15250 ( .A(n10256), .Y(n10251) );
  NOR2XL U15251 ( .A(n10254), .B(n10260), .Y(n10262) );
  INVXL U15252 ( .A(M2_U3_U1_enc_tree_4__4__16_), .Y(n10254) );
  OAI22XL U15253 ( .A0(n10247), .A1(n10272), .B0(M2_U3_U1_enc_tree_1__4__16_), 
        .B1(M2_U4_U1_enc_tree_1__4__16_), .Y(n10269) );
  NOR2XL U15254 ( .A(n10271), .B(n10270), .Y(n10247) );
  XOR2XL U15255 ( .A(n10267), .B(n10266), .Y(n10268) );
  NAND2XL U15256 ( .A(n10705), .B(n10704), .Y(n10272) );
  XOR2XL U15257 ( .A(n10271), .B(n10270), .Y(n10273) );
  INVXL U15258 ( .A(n10278), .Y(n10282) );
  XNOR2XL U15259 ( .A(n10705), .B(n10704), .Y(n10707) );
  INVX1 U15260 ( .A(n12688), .Y(n4940) );
  OAI22XL U15261 ( .A0(n12759), .A1(n12758), .B0(n12760), .B1(n12751), .Y(
        n12761) );
  OAI22XL U15262 ( .A0(n12535), .A1(M3_mult_x_15_b_21_), .B0(n12995), .B1(
        n3202), .Y(n12762) );
  NAND2XL U15263 ( .A(n12792), .B(n12791), .Y(n12822) );
  CMPR32X1 U15264 ( .A(n12710), .B(n12709), .C(n12708), .CO(n12725), .S(n12719) );
  OAI22XL U15265 ( .A0(n12715), .A1(n12699), .B0(n12746), .B1(n12714), .Y(
        n12710) );
  OAI2BB1XL U15266 ( .A0N(n12718), .A1N(n12717), .B0(n12716), .Y(n12726) );
  OAI22XL U15267 ( .A0(n12715), .A1(n12714), .B0(n12746), .B1(n12732), .Y(
        n12727) );
  OAI22XL U15268 ( .A0(n12759), .A1(n12729), .B0(n12760), .B1(n12745), .Y(
        n12744) );
  AOI21XL U15269 ( .A0(n13351), .A1(n13350), .B0(n13349), .Y(n13352) );
  OAI21XL U15270 ( .A0(n13346), .A1(n13345), .B0(n13344), .Y(n13351) );
  INVXL U15271 ( .A(n13664), .Y(n13604) );
  CLKINVX3 U15272 ( .A(n13661), .Y(n5286) );
  NOR2X2 U15273 ( .A(n14624), .B(n5280), .Y(n5150) );
  INVXL U15274 ( .A(n14370), .Y(n14374) );
  XNOR2XL U15275 ( .A(n14372), .B(n14371), .Y(n14373) );
  INVXL U15276 ( .A(n14376), .Y(n14381) );
  INVXL U15277 ( .A(n14377), .Y(n14380) );
  NAND2XL U15278 ( .A(n14479), .B(n14478), .Y(n14387) );
  XOR2XL U15279 ( .A(n14386), .B(n14385), .Y(n14388) );
  NAND2XL U15280 ( .A(n14376), .B(n14377), .Y(n14384) );
  XOR2XL U15281 ( .A(n14392), .B(n14391), .Y(n14393) );
  XOR2XL U15282 ( .A(n14390), .B(n14389), .Y(n14391) );
  INVXL U15283 ( .A(n24105), .Y(n14470) );
  INVXL U15284 ( .A(n14625), .Y(n14605) );
  NAND2XL U15285 ( .A(n17776), .B(n4885), .Y(n4650) );
  OR2XL U15286 ( .A(n17776), .B(n4885), .Y(n4883) );
  INVXL U15287 ( .A(n24376), .Y(n11618) );
  NAND2X1 U15288 ( .A(n6119), .B(n6118), .Y(n6117) );
  NAND2X1 U15289 ( .A(n5035), .B(n5034), .Y(n17653) );
  NAND2XL U15290 ( .A(n17599), .B(n17598), .Y(n5034) );
  ADDFX2 U15291 ( .A(n18602), .B(n18601), .CI(n18600), .CO(n18617), .S(n18612)
         );
  OAI22XL U15292 ( .A0(n18624), .A1(n18484), .B0(n18625), .B1(n18604), .Y(
        n18602) );
  NAND2X1 U15293 ( .A(n17645), .B(n6158), .Y(n6157) );
  OAI22XL U15294 ( .A0(n18721), .A1(M3_mult_x_15_b_21_), .B0(n17512), .B1(
        n3202), .Y(n18668) );
  OAI22XL U15295 ( .A0(n18659), .A1(n25883), .B0(n17832), .B1(n18658), .Y(
        n18667) );
  INVXL U15296 ( .A(n14509), .Y(n14510) );
  NAND2XL U15297 ( .A(n14341), .B(n14340), .Y(n14515) );
  NAND2XL U15298 ( .A(n14339), .B(n14338), .Y(n14509) );
  INVXL U15299 ( .A(n14506), .Y(n14511) );
  AOI2BB1XL U15300 ( .A0N(n20436), .A1N(n8955), .B0(n20435), .Y(n8956) );
  AOI2BB1XL U15301 ( .A0N(n8954), .A1N(n20440), .B0(n20439), .Y(n8955) );
  AOI2BB1XL U15302 ( .A0N(n8953), .A1N(n9015), .B0(n20443), .Y(n8954) );
  NAND2XL U15303 ( .A(n8765), .B(n8764), .Y(n8766) );
  INVXL U15304 ( .A(n8763), .Y(n8765) );
  AOI21XL U15305 ( .A0(n8860), .A1(n8859), .B0(n8858), .Y(n8861) );
  INVXL U15306 ( .A(n8854), .Y(n8857) );
  NAND2XL U15307 ( .A(n8853), .B(n8859), .Y(n8862) );
  INVX1 U15308 ( .A(n8783), .Y(n8863) );
  INVXL U15309 ( .A(n8875), .Y(n8838) );
  INVXL U15310 ( .A(n8876), .Y(n8877) );
  NAND2XL U15311 ( .A(n8875), .B(n8878), .Y(n8881) );
  AOI21XL U15312 ( .A0(n8825), .A1(n8823), .B0(n3155), .Y(n8824) );
  INVXL U15313 ( .A(n8830), .Y(n8872) );
  INVXL U15314 ( .A(n24063), .Y(n20143) );
  INVXL U15315 ( .A(n20204), .Y(n20140) );
  INVXL U15316 ( .A(n20203), .Y(n20206) );
  NAND2XL U15317 ( .A(n19867), .B(n19866), .Y(n19868) );
  INVXL U15318 ( .A(n19865), .Y(n19867) );
  NAND2XL U15319 ( .A(n19854), .B(n19853), .Y(n19855) );
  INVXL U15320 ( .A(n19852), .Y(n19854) );
  NAND2XL U15321 ( .A(n19880), .B(n19879), .Y(n19881) );
  INVXL U15322 ( .A(n19878), .Y(n19880) );
  NAND2XL U15323 ( .A(n19885), .B(n19884), .Y(n19886) );
  INVXL U15324 ( .A(n19883), .Y(n19885) );
  NAND2XL U15325 ( .A(n19858), .B(n19857), .Y(n19859) );
  NAND2XL U15326 ( .A(n19875), .B(n19874), .Y(n19876) );
  INVXL U15327 ( .A(n19870), .Y(n19873) );
  NOR2XL U15328 ( .A(n24986), .B(n20201), .Y(n20178) );
  NOR2XL U15329 ( .A(n3030), .B(n20176), .Y(n20179) );
  INVXL U15330 ( .A(n20196), .Y(n20176) );
  INVXL U15331 ( .A(n20195), .Y(n20198) );
  NOR2XL U15332 ( .A(n24986), .B(n20219), .Y(n20220) );
  NAND2XL U15333 ( .A(n20014), .B(n20013), .Y(n20015) );
  INVXL U15334 ( .A(n20012), .Y(n20014) );
  NAND2XL U15335 ( .A(n19995), .B(n19994), .Y(n19996) );
  INVXL U15336 ( .A(n19993), .Y(n19995) );
  INVXL U15337 ( .A(n24716), .Y(n24746) );
  NAND2XL U15338 ( .A(n19845), .B(n19984), .Y(n19846) );
  INVXL U15339 ( .A(n19985), .Y(n19845) );
  INVXL U15340 ( .A(n19959), .Y(n20001) );
  NOR2XL U15341 ( .A(n24986), .B(n20218), .Y(n20189) );
  INVXL U15342 ( .A(n20149), .Y(n20153) );
  NAND2XL U15343 ( .A(n25269), .B(n15761), .Y(n15756) );
  INVXL U15344 ( .A(n15835), .Y(n15838) );
  INVXL U15345 ( .A(n15836), .Y(n15753) );
  NAND2XL U15346 ( .A(n25269), .B(n15772), .Y(n15752) );
  NAND2XL U15347 ( .A(n25269), .B(n15835), .Y(n15805) );
  NOR2XL U15348 ( .A(n15772), .B(n15754), .Y(n15699) );
  NOR2XL U15349 ( .A(n15764), .B(n15830), .Y(n15802) );
  INVXL U15350 ( .A(n15861), .Y(n15800) );
  INVXL U15351 ( .A(n21000), .Y(n15911) );
  INVXL U15352 ( .A(n15626), .Y(n15627) );
  NAND2XL U15353 ( .A(n15625), .B(n15628), .Y(n15631) );
  NOR2XL U15354 ( .A(n15764), .B(n15831), .Y(n15832) );
  INVXL U15355 ( .A(n15761), .Y(n15767) );
  NAND2XL U15356 ( .A(n6216), .B(n22095), .Y(n22096) );
  NAND2XL U15357 ( .A(n22127), .B(n22126), .Y(n22129) );
  INVXL U15358 ( .A(n22302), .Y(n22236) );
  INVXL U15359 ( .A(n21625), .Y(n21791) );
  AOI2BB2XL U15360 ( .B0(n23116), .B1(n21870), .A0N(n21628), .A1N(n21871), .Y(
        n21714) );
  NAND2XL U15361 ( .A(n21628), .B(n21880), .Y(n21462) );
  AOI21XL U15362 ( .A0(n21783), .A1(n21560), .B0(n3037), .Y(n21710) );
  NOR2XL U15363 ( .A(n21582), .B(n21700), .Y(n21744) );
  AOI2BB2XL U15364 ( .B0(n23116), .B1(n21875), .A0N(n21628), .A1N(n21876), .Y(
        n21698) );
  AOI2BB2XL U15365 ( .B0(n23116), .B1(n21552), .A0N(n21628), .A1N(n21553), .Y(
        n21699) );
  INVXL U15366 ( .A(n21793), .Y(n21672) );
  NAND2XL U15367 ( .A(n3020), .B(n21961), .Y(n21515) );
  NAND2XL U15368 ( .A(n3020), .B(n21982), .Y(n21521) );
  AOI2BB2XL U15369 ( .B0(n23116), .B1(n21530), .A0N(n21628), .A1N(n21531), .Y(
        n21683) );
  NAND2XL U15370 ( .A(n21367), .B(n21434), .Y(n21368) );
  NAND2XL U15371 ( .A(n21372), .B(n21409), .Y(n21373) );
  NAND2XL U15372 ( .A(n21371), .B(n21405), .Y(n21374) );
  NAND2XL U15373 ( .A(n21356), .B(n21425), .Y(n21357) );
  NAND2XL U15374 ( .A(n21338), .B(n21517), .Y(n21339) );
  NAND2XL U15375 ( .A(n21343), .B(n21508), .Y(n21344) );
  NAND2XL U15376 ( .A(n21342), .B(n21520), .Y(n21345) );
  NAND2XL U15377 ( .A(n21351), .B(n21511), .Y(n21352) );
  INVXL U15378 ( .A(n15177), .Y(n15222) );
  NOR2XL U15379 ( .A(n15169), .B(n15154), .Y(n14783) );
  NAND2XL U15380 ( .A(n15665), .B(n15676), .Y(n15666) );
  NAND2XL U15381 ( .A(n15662), .B(n15675), .Y(n15663) );
  INVXL U15382 ( .A(n15676), .Y(n15661) );
  AOI21XL U15383 ( .A0(n15610), .A1(n15478), .B0(n15469), .Y(n15470) );
  INVXL U15384 ( .A(n15477), .Y(n15469) );
  NAND2XL U15385 ( .A(n15603), .B(n15478), .Y(n15471) );
  NAND2XL U15386 ( .A(n15455), .B(n15454), .Y(n15473) );
  NAND2XL U15387 ( .A(n15603), .B(n15601), .Y(n15457) );
  NAND2XL U15388 ( .A(n15464), .B(n15463), .Y(n15605) );
  INVXL U15389 ( .A(n22244), .Y(n22277) );
  INVXL U15390 ( .A(n22247), .Y(n22276) );
  INVXL U15391 ( .A(n22254), .Y(n22335) );
  NAND2XL U15392 ( .A(n22099), .B(n22112), .Y(n22100) );
  INVXL U15393 ( .A(n22113), .Y(n22098) );
  NAND2XL U15394 ( .A(n22102), .B(n22113), .Y(n22103) );
  NOR2X1 U15395 ( .A(n22213), .B(n22258), .Y(n22165) );
  AOI21XL U15396 ( .A0(n22013), .A1(n3222), .B0(n21849), .Y(n22012) );
  INVXL U15397 ( .A(n22018), .Y(n22060) );
  INVXL U15398 ( .A(n22130), .Y(n22132) );
  NOR2XL U15399 ( .A(n22207), .B(n22206), .Y(n22208) );
  NAND3XL U15400 ( .A(n22247), .B(n22295), .C(n22292), .Y(n22207) );
  NAND4XL U15401 ( .A(n22244), .B(n22205), .C(n22296), .D(n22297), .Y(n22206)
         );
  NOR2XL U15402 ( .A(n22204), .B(n22236), .Y(n22205) );
  NAND3XL U15403 ( .A(n22273), .B(n22286), .C(n22333), .Y(n22201) );
  AOI21XL U15404 ( .A0(n7920), .A1(n7919), .B0(n7918), .Y(n7955) );
  NAND2XL U15405 ( .A(n17137), .B(n17136), .Y(n17384) );
  INVXL U15406 ( .A(n10962), .Y(n10969) );
  INVXL U15407 ( .A(n10959), .Y(n11003) );
  INVXL U15408 ( .A(n23683), .Y(n7417) );
  INVXL U15409 ( .A(n23854), .Y(n7416) );
  INVXL U15410 ( .A(n10986), .Y(n10989) );
  INVXL U15411 ( .A(n10987), .Y(n10988) );
  INVXL U15412 ( .A(n10990), .Y(n11097) );
  INVXL U15413 ( .A(n11096), .Y(n10991) );
  NAND2XL U15414 ( .A(M6_mult_x_15_n500), .B(M6_mult_x_15_n508), .Y(n10993) );
  NOR2XL U15415 ( .A(M6_mult_x_15_n500), .B(M6_mult_x_15_n508), .Y(n10992) );
  NOR2XL U15416 ( .A(M6_mult_x_15_n518), .B(M6_mult_x_15_n527), .Y(n11031) );
  INVXL U15417 ( .A(n11028), .Y(n11346) );
  INVXL U15418 ( .A(n11345), .Y(n11029) );
  NAND2XL U15419 ( .A(M6_mult_x_15_n518), .B(M6_mult_x_15_n527), .Y(n11032) );
  XNOR2XL U15420 ( .A(n11099), .B(n11098), .Y(n20291) );
  NAND2XL U15421 ( .A(n11097), .B(n11096), .Y(n11098) );
  XNOR2XL U15422 ( .A(n11372), .B(n11037), .Y(n20290) );
  NAND2XL U15423 ( .A(n11356), .B(n11354), .Y(n11037) );
  AND2X2 U15424 ( .A(n4949), .B(n12901), .Y(n12918) );
  INVXL U15425 ( .A(n11036), .Y(n11356) );
  INVXL U15426 ( .A(n11354), .Y(n11355) );
  INVXL U15427 ( .A(n11006), .Y(n10952) );
  INVXL U15428 ( .A(n11021), .Y(n10951) );
  NAND2XL U15429 ( .A(M6_mult_x_15_n463), .B(M6_mult_x_15_n468), .Y(n10979) );
  NAND2XL U15430 ( .A(M6_mult_x_15_n462), .B(M6_mult_x_15_n457), .Y(n10974) );
  INVXL U15431 ( .A(n7768), .Y(n7770) );
  NAND2XL U15432 ( .A(M6_mult_x_15_n451), .B(M6_mult_x_15_n456), .Y(n10968) );
  NAND2XL U15433 ( .A(M6_mult_x_15_n450), .B(M6_mult_x_15_n446), .Y(n10964) );
  NOR2XL U15434 ( .A(M6_mult_x_15_n451), .B(M6_mult_x_15_n456), .Y(n10962) );
  INVXL U15435 ( .A(n11038), .Y(n11041) );
  INVXL U15436 ( .A(n11039), .Y(n11040) );
  INVXL U15437 ( .A(n11042), .Y(n11338) );
  INVXL U15438 ( .A(n11336), .Y(n11337) );
  NAND2XL U15439 ( .A(M6_mult_x_15_n538), .B(M6_mult_x_15_n548), .Y(n11341) );
  NOR2XL U15440 ( .A(M6_mult_x_15_n538), .B(M6_mult_x_15_n548), .Y(n11340) );
  XOR2XL U15441 ( .A(n11348), .B(n11347), .Y(n11468) );
  NAND2XL U15442 ( .A(n11346), .B(n11345), .Y(n11347) );
  XOR2XL U15443 ( .A(n11118), .B(n11117), .Y(n11466) );
  NAND2XL U15444 ( .A(n11116), .B(n11115), .Y(n11117) );
  INVXL U15445 ( .A(n11114), .Y(n11116) );
  NAND2XL U15446 ( .A(M6_mult_x_15_n469), .B(M6_mult_x_15_n475), .Y(n10999) );
  XNOR2XL U15447 ( .A(n11353), .B(n11352), .Y(n20289) );
  NAND2XL U15448 ( .A(n11351), .B(n11350), .Y(n11352) );
  AOI21XL U15449 ( .A0(n10936), .A1(n10935), .B0(n10934), .Y(n11106) );
  NOR2XL U15450 ( .A(n10933), .B(n10744), .Y(n10936) );
  XOR2XL U15451 ( .A(n22622), .B(n3221), .Y(M6_mult_x_15_n1194) );
  XNOR2XL U15452 ( .A(n11279), .B(n11278), .Y(n11332) );
  NAND2XL U15453 ( .A(n11277), .B(n11276), .Y(n11278) );
  OAI2BB1XL U15454 ( .A0N(n11263), .A1N(n11262), .B0(n11261), .Y(n11456) );
  NAND3XL U15455 ( .A(n11260), .B(n11264), .C(n11259), .Y(n11261) );
  AND2XL U15456 ( .A(n11272), .B(n11271), .Y(n11273) );
  NAND2X1 U15457 ( .A(n5612), .B(n5611), .Y(n6900) );
  NAND2XL U15458 ( .A(n6894), .B(n6895), .Y(n5611) );
  NOR2X1 U15459 ( .A(n5684), .B(n17389), .Y(n5683) );
  NOR2X1 U15460 ( .A(n17375), .B(n17387), .Y(n5684) );
  INVXL U15461 ( .A(n17387), .Y(n17390) );
  INVXL U15462 ( .A(n25162), .Y(n17198) );
  NAND2X1 U15463 ( .A(n16954), .B(n16955), .Y(n5829) );
  NOR2X1 U15464 ( .A(n16954), .B(n16955), .Y(n5831) );
  AOI21XL U15465 ( .A0(n10734), .A1(n10733), .B0(n10732), .Y(n10735) );
  XOR2XL U15466 ( .A(n10731), .B(n10730), .Y(n10733) );
  NAND2XL U15467 ( .A(n12959), .B(n12958), .Y(n13032) );
  AOI22XL U15468 ( .A0(n12957), .A1(n12956), .B0(n12955), .B1(n18810), .Y(
        n12958) );
  NAND2XL U15469 ( .A(n12960), .B(n12952), .Y(n12959) );
  INVXL U15470 ( .A(n12954), .Y(n12956) );
  NOR2XL U15471 ( .A(n12970), .B(n12969), .Y(n13034) );
  NAND2XL U15472 ( .A(n12968), .B(n12967), .Y(n12969) );
  INVXL U15473 ( .A(n12960), .Y(n12970) );
  XOR2XL U15474 ( .A(n12966), .B(n12965), .Y(n12967) );
  XOR2XL U15475 ( .A(n18840), .B(n13031), .Y(n13033) );
  NAND2XL U15476 ( .A(n11362), .B(n11367), .Y(n11370) );
  NOR2XL U15477 ( .A(M6_mult_x_15_n560), .B(M6_mult_x_15_n570), .Y(n11101) );
  NAND2XL U15478 ( .A(M6_mult_x_15_n571), .B(M6_mult_x_15_n581), .Y(n11115) );
  NOR2XL U15479 ( .A(M6_mult_x_15_n571), .B(M6_mult_x_15_n581), .Y(n11114) );
  NAND2XL U15480 ( .A(M6_mult_x_15_n560), .B(M6_mult_x_15_n570), .Y(n11102) );
  INVXL U15481 ( .A(n10983), .Y(n11118) );
  XNOR2XL U15482 ( .A(n11339), .B(n11043), .Y(n11465) );
  NAND2XL U15483 ( .A(n11338), .B(n11336), .Y(n11043) );
  INVXL U15484 ( .A(M5_U3_U1_enc_tree_0__4__16_), .Y(n17414) );
  INVXL U15485 ( .A(M5_U3_U1_enc_tree_0__2__12_), .Y(
        M5_U3_U1_enc_tree_0__3__8_) );
  AOI21XL U15486 ( .A0(n4888), .A1(n3210), .B0(M4_a_12_), .Y(
        M4_U3_U1_enc_tree_0__1__18_) );
  AOI21XL U15487 ( .A0(n18658), .A1(n5471), .B0(M4_a_20_), .Y(
        M4_U3_U1_enc_tree_0__1__10_) );
  OR2XL U15488 ( .A(M4_U3_U1_or2_tree_0__2__16_), .B(
        M4_U3_U1_or2_tree_0__2__24_), .Y(n26154) );
  INVXL U15489 ( .A(M3_U4_U1_or2_tree_0__2__24_), .Y(M3_U4_U1_or2_inv_0__24_)
         );
  AND2XL U15490 ( .A(M4_U3_U1_enc_tree_3__3__16_), .B(
        M4_U3_U1_enc_tree_3__3__24_), .Y(n18811) );
  NOR2XL U15491 ( .A(n18810), .B(n18811), .Y(n18809) );
  XOR2XL U15492 ( .A(n18806), .B(n18805), .Y(n18807) );
  INVXL U15493 ( .A(n18802), .Y(n18806) );
  INVXL U15494 ( .A(n18808), .Y(n18813) );
  NAND2XL U15495 ( .A(n18840), .B(n18839), .Y(n18823) );
  NAND2XL U15496 ( .A(n18808), .B(n18809), .Y(n18816) );
  XOR2XL U15497 ( .A(n18820), .B(n18819), .Y(n18826) );
  XOR2XL U15498 ( .A(n18818), .B(n18817), .Y(n18819) );
  INVXL U15499 ( .A(n11044), .Y(n11362) );
  NAND2XL U15500 ( .A(M6_mult_x_15_n438), .B(M6_mult_x_15_n441), .Y(n11009) );
  NOR2XL U15501 ( .A(M6_mult_x_15_n445), .B(M6_mult_x_15_n442), .Y(n10959) );
  INVXL U15502 ( .A(n11004), .Y(n10956) );
  INVXL U15503 ( .A(n11015), .Y(n10955) );
  NAND2XL U15504 ( .A(n11121), .B(n11120), .Y(n11122) );
  INVXL U15505 ( .A(n11119), .Y(n11121) );
  AOI31XL U15506 ( .A0(n11457), .A1(n20957), .A2(n11456), .B0(n11455), .Y(
        n11458) );
  INVXL U15507 ( .A(n11454), .Y(n11457) );
  AOI211XL U15508 ( .A0(n11453), .A1(n11452), .B0(n11451), .C0(n11450), .Y(
        n11454) );
  INVXL U15509 ( .A(n11092), .Y(n11375) );
  AOI21XL U15510 ( .A0(n23150), .A1(n11071), .B0(n23093), .Y(n11091) );
  XOR2XL U15511 ( .A(n22523), .B(n3119), .Y(M6_mult_x_15_n1029) );
  INVXL U15512 ( .A(n23096), .Y(M6_mult_x_15_n1006) );
  INVXL U15513 ( .A(n23077), .Y(M6_mult_x_15_n1005) );
  AOI21XL U15514 ( .A0(n23150), .A1(n3218), .B0(n23074), .Y(n23075) );
  AOI21XL U15515 ( .A0(n11024), .A1(n11023), .B0(n11022), .Y(n11371) );
  NAND2XL U15516 ( .A(n11007), .B(n11024), .Y(n11363) );
  INVXL U15517 ( .A(n11374), .Y(n11394) );
  INVXL U15518 ( .A(n23150), .Y(n11373) );
  INVXL U15519 ( .A(n11387), .Y(n11388) );
  NOR3XL U15520 ( .A(n23678), .B(n25835), .C(n11331), .Y(n6218) );
  NAND3BXL U15521 ( .AN(n24443), .B(n11330), .C(n11405), .Y(n11331) );
  INVXL U15522 ( .A(n20457), .Y(n20460) );
  INVXL U15523 ( .A(n20453), .Y(n20456) );
  NAND2XL U15524 ( .A(n3067), .B(n20454), .Y(n20455) );
  INVXL U15525 ( .A(n20543), .Y(n20399) );
  NAND2XL U15526 ( .A(n3067), .B(n20449), .Y(n20398) );
  NAND2XL U15527 ( .A(n14427), .B(y10[28]), .Y(n9132) );
  NOR2XL U15528 ( .A(n3124), .B(n20463), .Y(n20416) );
  INVXL U15529 ( .A(n20458), .Y(n20414) );
  INVXL U15530 ( .A(n20400), .Y(n20580) );
  NAND2XL U15531 ( .A(n7741), .B(n7790), .Y(n7742) );
  INVXL U15532 ( .A(n7791), .Y(n7741) );
  INVXL U15533 ( .A(n7724), .Y(n7702) );
  NAND2XL U15534 ( .A(n7717), .B(n7716), .Y(n7723) );
  INVXL U15535 ( .A(n10521), .Y(n10638) );
  AOI21XL U15536 ( .A0(n10233), .A1(n10224), .B0(n10183), .Y(n10184) );
  NAND2XL U15537 ( .A(n10553), .B(n10552), .Y(n10645) );
  OR2X2 U15538 ( .A(n10643), .B(n10656), .Y(n5248) );
  NOR2XL U15539 ( .A(n10581), .B(n10656), .Y(n5007) );
  NAND2XL U15540 ( .A(n10596), .B(n10601), .Y(n10581) );
  INVXL U15541 ( .A(n10600), .Y(n10579) );
  NAND2XL U15542 ( .A(n10560), .B(n10559), .Y(n10583) );
  NAND2XL U15543 ( .A(n10593), .B(n10592), .Y(n10594) );
  INVXL U15544 ( .A(n10591), .Y(n10593) );
  NAND2X1 U15545 ( .A(n11920), .B(n4974), .Y(n4972) );
  INVX1 U15546 ( .A(n12979), .Y(n12859) );
  INVX1 U15547 ( .A(n12890), .Y(n12914) );
  NAND2X1 U15548 ( .A(n12853), .B(n12611), .Y(n12839) );
  XNOR2X1 U15549 ( .A(n12705), .B(n12707), .Y(n6001) );
  INVX1 U15550 ( .A(n12995), .Y(n12994) );
  INVX1 U15551 ( .A(n12978), .Y(n12834) );
  INVXL U15552 ( .A(n12829), .Y(n12831) );
  XNOR2X1 U15553 ( .A(n14558), .B(n14557), .Y(n14669) );
  NAND2XL U15554 ( .A(n14550), .B(n14570), .Y(n14554) );
  INVXL U15555 ( .A(n24110), .Y(n18788) );
  NAND2XL U15556 ( .A(n14360), .B(n14359), .Y(n14361) );
  NAND2X2 U15557 ( .A(n14309), .B(n14310), .Y(n14591) );
  INVXL U15558 ( .A(n18942), .Y(n18955) );
  NAND2XL U15559 ( .A(n14328), .B(n14327), .Y(n14538) );
  INVX1 U15560 ( .A(n17229), .Y(n5713) );
  INVXL U15561 ( .A(n19003), .Y(n18985) );
  NAND2XL U15562 ( .A(n18707), .B(n18706), .Y(n18989) );
  INVXL U15563 ( .A(n14618), .Y(n14620) );
  NAND2XL U15564 ( .A(n14651), .B(n14650), .Y(n14652) );
  NOR2XL U15565 ( .A(n9016), .B(n9028), .Y(n8947) );
  NAND4XL U15566 ( .A(n20562), .B(n20458), .C(n20542), .D(n20453), .Y(n9025)
         );
  NOR2XL U15567 ( .A(n20156), .B(n24063), .Y(n20077) );
  INVXL U15568 ( .A(n24889), .Y(n24851) );
  INVXL U15569 ( .A(n24938), .Y(n24891) );
  NAND2XL U15570 ( .A(n3030), .B(n24889), .Y(n24890) );
  NOR2XL U15571 ( .A(n3030), .B(n24985), .Y(n24988) );
  INVXL U15572 ( .A(n25344), .Y(n24985) );
  INVXL U15573 ( .A(n15826), .Y(n15829) );
  NAND2XL U15574 ( .A(n25269), .B(n15827), .Y(n15828) );
  INVXL U15575 ( .A(n15860), .Y(n15863) );
  INVXL U15576 ( .A(n15923), .Y(n15797) );
  INVXL U15577 ( .A(n15920), .Y(n15921) );
  INVXL U15578 ( .A(n22202), .Y(n22307) );
  NAND2XL U15579 ( .A(n22090), .B(n22089), .Y(n22091) );
  NAND2XL U15580 ( .A(n22188), .B(n22198), .Y(n22187) );
  NOR2XL U15581 ( .A(n21366), .B(n21430), .Y(n21325) );
  AOI21XL U15582 ( .A0(n14769), .A1(n14768), .B0(n14767), .Y(n14792) );
  OAI22XL U15583 ( .A0(n22343), .A1(n22318), .B0(n22317), .B1(n3129), .Y(
        n22367) );
  NOR2XL U15584 ( .A(n22337), .B(n22336), .Y(n22427) );
  NOR2XL U15585 ( .A(n22308), .B(n22335), .Y(n22336) );
  INVXL U15586 ( .A(n22333), .Y(n22334) );
  AOI21XL U15587 ( .A0(n22338), .A1(n3129), .B0(n22290), .Y(n22420) );
  NOR2XL U15588 ( .A(n22318), .B(n3129), .Y(n22319) );
  INVXL U15589 ( .A(n22448), .Y(n22449) );
  INVXL U15590 ( .A(n22256), .Y(n22450) );
  NAND2XL U15591 ( .A(n21331), .B(w1[23]), .Y(n21305) );
  AOI2BB1XL U15592 ( .A0N(n22145), .A1N(n22244), .B0(n22247), .Y(n22146) );
  NAND2XL U15593 ( .A(n22032), .B(n22031), .Y(n22033) );
  INVXL U15594 ( .A(n22030), .Y(n22032) );
  NAND2XL U15595 ( .A(n22066), .B(n22064), .Y(n22028) );
  INVXL U15596 ( .A(n22063), .Y(n22026) );
  NAND2XL U15597 ( .A(n22037), .B(n22036), .Y(n22038) );
  INVXL U15598 ( .A(n22035), .Y(n22037) );
  NAND2XL U15599 ( .A(n22054), .B(n22053), .Y(n22055) );
  INVXL U15600 ( .A(n22052), .Y(n22054) );
  NAND2XL U15601 ( .A(n22073), .B(n22072), .Y(n22074) );
  INVXL U15602 ( .A(n22071), .Y(n22073) );
  NOR4XL U15603 ( .A(n23404), .B(n23400), .C(n23408), .D(n23416), .Y(n22182)
         );
  NAND3XL U15604 ( .A(n22448), .B(n22272), .C(n22254), .Y(n22210) );
  NAND4XL U15605 ( .A(n22208), .B(n22287), .C(n22285), .D(n22282), .Y(n22209)
         );
  XOR2XL U15606 ( .A(n9159), .B(n10674), .Y(n9161) );
  XNOR2XL U15607 ( .A(n10982), .B(n10981), .Y(n20288) );
  NAND2XL U15608 ( .A(n10980), .B(n10979), .Y(n10981) );
  INVXL U15609 ( .A(n10978), .Y(n10980) );
  XNOR2XL U15610 ( .A(n10971), .B(n10970), .Y(n20287) );
  NAND2XL U15611 ( .A(n10969), .B(n10968), .Y(n10970) );
  NAND2XL U15612 ( .A(n11003), .B(n11008), .Y(n10960) );
  NAND2XL U15613 ( .A(n5604), .B(w2[30]), .Y(n7386) );
  NAND2XL U15614 ( .A(n7389), .B(y10[30]), .Y(n7385) );
  NAND2XL U15615 ( .A(n9119), .B(n14407), .Y(n9120) );
  NAND2XL U15616 ( .A(n25233), .B(sigma10[24]), .Y(n9119) );
  NAND2XL U15617 ( .A(n9126), .B(n14410), .Y(n9127) );
  NAND2XL U15618 ( .A(n25233), .B(sigma10[26]), .Y(n9126) );
  NAND2XL U15619 ( .A(n9111), .B(n14416), .Y(n9112) );
  NAND2XL U15620 ( .A(n25233), .B(sigma10[30]), .Y(n9111) );
  NAND2XL U15621 ( .A(n4856), .B(target_temp[27]), .Y(n14440) );
  NAND2XL U15622 ( .A(n4826), .B(target_temp[28]), .Y(n14436) );
  NAND2XL U15623 ( .A(n21166), .B(sigma10[30]), .Y(n11552) );
  INVXL U15624 ( .A(n17316), .Y(n17318) );
  NOR2XL U15625 ( .A(n20293), .B(n20292), .Y(n23914) );
  XOR2XL U15626 ( .A(n11035), .B(n11034), .Y(n23916) );
  NAND2XL U15627 ( .A(n11033), .B(n11032), .Y(n11034) );
  AOI21XL U15628 ( .A0(n11030), .A1(n11346), .B0(n11029), .Y(n11035) );
  INVXL U15629 ( .A(n11031), .Y(n11033) );
  NAND2XL U15630 ( .A(n23916), .B(n23914), .Y(n23501) );
  INVXL U15631 ( .A(n20291), .Y(n23503) );
  NAND2XL U15632 ( .A(n23498), .B(n23497), .Y(n23903) );
  INVXL U15633 ( .A(n20290), .Y(n23905) );
  INVXL U15634 ( .A(n20288), .Y(n20771) );
  NAND2X1 U15635 ( .A(n12918), .B(n12914), .Y(n12921) );
  NOR2XL U15636 ( .A(n23905), .B(n23903), .Y(n23598) );
  XOR2XL U15637 ( .A(n11361), .B(n11360), .Y(n23599) );
  NAND2XL U15638 ( .A(n11359), .B(n11358), .Y(n11360) );
  INVXL U15639 ( .A(n11357), .Y(n11359) );
  NAND2XL U15640 ( .A(n20766), .B(n20765), .Y(n20820) );
  INVXL U15641 ( .A(n20287), .Y(n20822) );
  INVXL U15642 ( .A(n7746), .Y(n7744) );
  NAND2XL U15643 ( .A(n10965), .B(n10964), .Y(n10966) );
  NAND2XL U15644 ( .A(n23541), .B(n23540), .Y(n20296) );
  INVXL U15645 ( .A(n20286), .Y(n20298) );
  NAND2XL U15646 ( .A(n7805), .B(n7807), .Y(n7810) );
  NOR2XL U15647 ( .A(n23465), .B(n23463), .Y(n11472) );
  XOR2XL U15648 ( .A(n11344), .B(n11343), .Y(n11473) );
  NAND2XL U15649 ( .A(n11342), .B(n11341), .Y(n11343) );
  AOI21XL U15650 ( .A0(n11339), .A1(n11338), .B0(n11337), .Y(n11344) );
  INVXL U15651 ( .A(n11340), .Y(n11342) );
  NAND2XL U15652 ( .A(n11473), .B(n11472), .Y(n20292) );
  INVXL U15653 ( .A(n11468), .Y(n20293) );
  XNOR2XL U15654 ( .A(n11113), .B(n11112), .Y(n19080) );
  NAND2XL U15655 ( .A(n11111), .B(n11110), .Y(n11112) );
  INVXL U15656 ( .A(n11109), .Y(n11111) );
  INVXL U15657 ( .A(n11466), .Y(n19081) );
  NOR2XL U15658 ( .A(n23596), .B(n23594), .Y(n23895) );
  XNOR2XL U15659 ( .A(n11002), .B(n11001), .Y(n23896) );
  NAND2XL U15660 ( .A(n11000), .B(n10999), .Y(n11001) );
  NAND2XL U15661 ( .A(n23599), .B(n23598), .Y(n23594) );
  INVXL U15662 ( .A(n20289), .Y(n23596) );
  NOR2XL U15663 ( .A(M6_mult_x_15_n604), .B(M6_mult_x_15_n614), .Y(n11126) );
  INVXL U15664 ( .A(n11106), .Y(n11279) );
  INVXL U15665 ( .A(n11124), .Y(n11277) );
  INVXL U15666 ( .A(n11276), .Y(n11125) );
  NAND2XL U15667 ( .A(M6_mult_x_15_n604), .B(M6_mult_x_15_n614), .Y(n11127) );
  AOI21XL U15668 ( .A0(n11335), .A1(n11334), .B0(n11333), .Y(n11459) );
  NAND2XL U15669 ( .A(n11456), .B(n11451), .Y(n11335) );
  NOR2XL U15670 ( .A(n11332), .B(n6218), .Y(n11333) );
  INVXL U15671 ( .A(n20957), .Y(n11334) );
  NOR2XL U15672 ( .A(n17203), .B(n25222), .Y(n17202) );
  INVXL U15673 ( .A(n19080), .Y(n19063) );
  NOR2X2 U15674 ( .A(n17120), .B(n17119), .Y(n17348) );
  NAND2XL U15675 ( .A(n11377), .B(n11376), .Y(n11387) );
  NAND2XL U15676 ( .A(n23468), .B(n23467), .Y(n23463) );
  INVXL U15677 ( .A(n11465), .Y(n23465) );
  NAND2XL U15678 ( .A(n17151), .B(n17150), .Y(n17152) );
  NAND2XL U15679 ( .A(n11463), .B(n11462), .Y(n19065) );
  NOR2XL U15680 ( .A(n11463), .B(n11462), .Y(n19064) );
  NOR2XL U15681 ( .A(M6_mult_x_15_n437), .B(M6_mult_x_15_n435), .Y(n11044) );
  NAND2XL U15682 ( .A(M6_mult_x_15_n434), .B(n11093), .Y(n11365) );
  NAND2XL U15683 ( .A(M6_mult_x_15_n437), .B(M6_mult_x_15_n435), .Y(n11364) );
  XOR2XL U15684 ( .A(n11396), .B(n11395), .Y(n11397) );
  NAND2XL U15685 ( .A(n11386), .B(n11389), .Y(n11392) );
  AOI2BB1X1 U15686 ( .A0N(n17241), .A1N(n17242), .B0(n17240), .Y(n17243) );
  NAND2XL U15687 ( .A(n21166), .B(sigma10[28]), .Y(n11570) );
  NAND2XL U15688 ( .A(n21166), .B(sigma10[24]), .Y(n11558) );
  NAND2XL U15689 ( .A(n3071), .B(n20592), .Y(n20593) );
  AOI2BB2XL U15690 ( .B0(n20505), .B1(n20473), .A0N(n20555), .A1N(n20473), .Y(
        n20426) );
  NOR2XL U15691 ( .A(n20408), .B(n20597), .Y(n20409) );
  NOR2XL U15692 ( .A(n20406), .B(n20405), .Y(n20407) );
  NOR2XL U15693 ( .A(n3124), .B(n20579), .Y(n20405) );
  NAND2XL U15694 ( .A(n19564), .B(n19319), .Y(n19320) );
  INVXL U15695 ( .A(n19310), .Y(n19313) );
  INVXL U15696 ( .A(n19314), .Y(n19317) );
  NAND2XL U15697 ( .A(n3041), .B(n19315), .Y(n19316) );
  NAND2XL U15698 ( .A(n19564), .B(n19323), .Y(n19324) );
  NAND2X1 U15699 ( .A(n20502), .B(n20576), .Y(n20538) );
  NAND2XL U15700 ( .A(n5604), .B(w2[26]), .Y(n7377) );
  NAND2XL U15701 ( .A(n6733), .B(y10[26]), .Y(n7376) );
  NAND2XL U15702 ( .A(n6733), .B(y10[28]), .Y(n7380) );
  NAND2XL U15703 ( .A(n5604), .B(w2[28]), .Y(n7381) );
  NAND2XL U15704 ( .A(n20988), .B(n19074), .Y(n5316) );
  NAND2X1 U15705 ( .A(n23495), .B(n20988), .Y(n5320) );
  NAND2X1 U15706 ( .A(n23489), .B(n19098), .Y(n19100) );
  NAND2XL U15707 ( .A(n19074), .B(n19073), .Y(n20990) );
  NOR2XL U15708 ( .A(n25267), .B(n3070), .Y(n25275) );
  NAND2XL U15709 ( .A(n25271), .B(n25270), .Y(n25272) );
  NOR2XL U15710 ( .A(n25266), .B(n3125), .Y(n25277) );
  INVXL U15711 ( .A(n25268), .Y(n15784) );
  AND2XL U15712 ( .A(n10706), .B(n10708), .Y(n4690) );
  NAND2X1 U15713 ( .A(n5281), .B(n5247), .Y(n5075) );
  NAND2X2 U15714 ( .A(n20324), .B(n20321), .Y(n20966) );
  NOR2X1 U15715 ( .A(n12839), .B(n12834), .Y(n12845) );
  INVX1 U15716 ( .A(n12873), .Y(n6134) );
  NOR2XL U15717 ( .A(n12985), .B(n12866), .Y(n12973) );
  AOI21XL U15718 ( .A0(n18935), .A1(n3000), .B0(n18934), .Y(n18936) );
  NOR2XL U15719 ( .A(n14480), .B(n14482), .Y(n14475) );
  INVXL U15720 ( .A(n20327), .Y(n20328) );
  NOR2XL U15721 ( .A(n18971), .B(n20658), .Y(n18970) );
  NAND2X1 U15722 ( .A(n18416), .B(n18417), .Y(n18882) );
  INVXL U15723 ( .A(n20975), .Y(n23444) );
  INVXL U15724 ( .A(n18870), .Y(n18873) );
  NAND2X1 U15725 ( .A(n20975), .B(n23447), .Y(n5275) );
  NOR2XL U15726 ( .A(n11623), .B(n25806), .Y(n11622) );
  AOI21X1 U15727 ( .A0(n14476), .A1(n5272), .B0(n5093), .Y(n5092) );
  INVXL U15728 ( .A(n14639), .Y(n14641) );
  INVX1 U15729 ( .A(n20661), .Y(n23707) );
  INVXL U15730 ( .A(n19015), .Y(n19017) );
  XNOR2X1 U15731 ( .A(n14681), .B(n14680), .Y(n23745) );
  NAND2XL U15732 ( .A(n14679), .B(n14678), .Y(n14680) );
  NOR2X1 U15733 ( .A(n3134), .B(n5388), .Y(n5384) );
  INVX1 U15734 ( .A(n23742), .Y(n5388) );
  INVXL U15735 ( .A(n14682), .Y(n23742) );
  INVXL U15736 ( .A(n20654), .Y(n20656) );
  NOR2BXL U15737 ( .AN(n24028), .B(n24027), .Y(n24033) );
  OAI22XL U15738 ( .A0(n20229), .A1(n3069), .B0(n20251), .B1(n20182), .Y(
        n24721) );
  NOR2XL U15739 ( .A(n25342), .B(n3032), .Y(n25347) );
  AND3XL U15740 ( .A(n25346), .B(n3032), .C(n25345), .Y(n6177) );
  NOR2XL U15741 ( .A(n25341), .B(n3069), .Y(n25349) );
  AOI2BB2XL U15742 ( .B0(n15893), .B1(n15745), .A0N(n15892), .A1N(n3125), .Y(
        n15928) );
  INVX1 U15743 ( .A(n23960), .Y(n15794) );
  AOI21XL U15744 ( .A0(n24921), .A1(n24920), .B0(n15688), .Y(n24922) );
  NAND2XL U15745 ( .A(n24919), .B(n3127), .Y(n24920) );
  INVXL U15746 ( .A(n24918), .Y(n24919) );
  NOR2XL U15747 ( .A(n25267), .B(n3127), .Y(n24966) );
  NAND2XL U15748 ( .A(n25010), .B(n25009), .Y(n25013) );
  NAND2XL U15749 ( .A(n25011), .B(n3127), .Y(n25012) );
  NAND2XL U15750 ( .A(n25269), .B(n25007), .Y(n25010) );
  INVXL U15751 ( .A(n22398), .Y(n22403) );
  NAND2XL U15752 ( .A(n22351), .B(n3079), .Y(n22345) );
  AOI21XL U15753 ( .A0(n21739), .A1(n21738), .B0(n21737), .Y(n22195) );
  NOR2XL U15754 ( .A(n22436), .B(n3129), .Y(n22261) );
  NOR2XL U15755 ( .A(n22411), .B(n3079), .Y(n22263) );
  INVXL U15756 ( .A(n21413), .Y(n21416) );
  NAND2XL U15757 ( .A(n23116), .B(n21414), .Y(n21415) );
  INVXL U15758 ( .A(n21430), .Y(n21433) );
  INVXL U15759 ( .A(n21434), .Y(n21437) );
  INVXL U15760 ( .A(n21425), .Y(n21428) );
  INVXL U15761 ( .A(n21405), .Y(n21408) );
  NAND2XL U15762 ( .A(n23116), .B(n21406), .Y(n21407) );
  OAI21XL U15763 ( .A0(n21519), .A1(n21412), .B0(n21411), .Y(n23120) );
  INVXL U15764 ( .A(n21409), .Y(n21412) );
  NAND2XL U15765 ( .A(n21628), .B(n21410), .Y(n21411) );
  NAND2XL U15766 ( .A(n21519), .B(n21418), .Y(n21419) );
  INVXL U15767 ( .A(n15730), .Y(n15731) );
  NAND2XL U15768 ( .A(n15729), .B(n15728), .Y(n15733) );
  OAI31XL U15769 ( .A0(n15920), .A1(n15923), .A2(n15727), .B0(n15726), .Y(
        n15728) );
  OAI21XL U15770 ( .A0(n15558), .A1(n14937), .B0(n14936), .Y(n23158) );
  NAND2XL U15771 ( .A(n15558), .B(n14935), .Y(n14936) );
  INVXL U15772 ( .A(n14926), .Y(n14929) );
  INVXL U15773 ( .A(n14930), .Y(n14933) );
  NAND2XL U15774 ( .A(n15190), .B(n14931), .Y(n14932) );
  NAND2XL U15775 ( .A(n15190), .B(n14939), .Y(n14940) );
  INVXL U15776 ( .A(n14950), .Y(n14953) );
  INVXL U15777 ( .A(n14954), .Y(n14957) );
  INVXL U15778 ( .A(n14942), .Y(n14945) );
  OAI21X1 U15779 ( .A0(n15558), .A1(n14949), .B0(n14948), .Y(n23164) );
  NAND2XL U15780 ( .A(n15190), .B(n14947), .Y(n14948) );
  OAI21XL U15781 ( .A0(n15558), .A1(n14915), .B0(n14914), .Y(n24060) );
  NAND2XL U15782 ( .A(n22370), .B(n3130), .Y(n22371) );
  NAND2XL U15783 ( .A(n22359), .B(n3130), .Y(n22360) );
  NAND2XL U15784 ( .A(n22354), .B(n3130), .Y(n22355) );
  OAI22XL U15785 ( .A0(n3130), .A1(n22367), .B0(n22406), .B1(n3079), .Y(n22267) );
  NAND2XL U15786 ( .A(n22368), .B(n3130), .Y(n22251) );
  NOR2X1 U15787 ( .A(n22381), .B(n22124), .Y(n22271) );
  NAND2XL U15788 ( .A(n3079), .B(n22420), .Y(n22291) );
  NAND2XL U15789 ( .A(n22384), .B(n22124), .Y(n22312) );
  NAND2XL U15790 ( .A(n22324), .B(n22426), .Y(n22325) );
  NOR2BXL U15791 ( .AN(n22354), .B(n3130), .Y(n22386) );
  INVXL U15792 ( .A(n23337), .Y(n23330) );
  AOI2BB1XL U15793 ( .A0N(n22411), .A1N(n3130), .B0(n22124), .Y(n22412) );
  OAI22XL U15794 ( .A0(n22406), .A1(n3130), .B0(n3079), .B1(n22402), .Y(n22410) );
  NAND2BXL U15795 ( .AN(n22124), .B(n23113), .Y(n22418) );
  NAND2XL U15796 ( .A(n22427), .B(n22426), .Y(n22428) );
  NAND2XL U15797 ( .A(n22420), .B(n3130), .Y(n22431) );
  NAND2XL U15798 ( .A(n22373), .B(n3130), .Y(n22374) );
  NOR2XL U15799 ( .A(n22437), .B(n3129), .Y(n22438) );
  NOR2XL U15800 ( .A(n22436), .B(n22343), .Y(n22439) );
  NOR2XL U15801 ( .A(n22440), .B(n3079), .Y(n22441) );
  NAND2XL U15802 ( .A(n23341), .B(n23311), .Y(n23329) );
  NAND2XL U15803 ( .A(n22455), .B(n3130), .Y(n22456) );
  AOI21XL U15804 ( .A0(n22250), .A1(n22454), .B0(n22453), .Y(n22457) );
  NOR2XL U15805 ( .A(n22452), .B(n22451), .Y(n22453) );
  NOR2XL U15806 ( .A(n22308), .B(n22450), .Y(n22451) );
  NOR2XL U15807 ( .A(n3126), .B(n22449), .Y(n22452) );
  NAND2XL U15808 ( .A(n22351), .B(n3130), .Y(n22352) );
  NAND2XL U15809 ( .A(n21331), .B(temp0[23]), .Y(n21306) );
  INVXL U15810 ( .A(n21417), .Y(n21420) );
  INVXL U15811 ( .A(n8207), .Y(n8210) );
  NAND2XL U15812 ( .A(n3040), .B(n8189), .Y(n8190) );
  NAND2XL U15813 ( .A(n8482), .B(n8193), .Y(n8194) );
  INVXL U15814 ( .A(n8199), .Y(n8202) );
  INVXL U15815 ( .A(n8195), .Y(n8198) );
  INVXL U15816 ( .A(n8180), .Y(n8183) );
  INVXL U15817 ( .A(n8184), .Y(n8187) );
  NAND2XL U15818 ( .A(n3111), .B(sigma10[23]), .Y(n11602) );
  NOR4BXL U15819 ( .AN(n20288), .B(n11383), .C(n11382), .D(n11381), .Y(n11384)
         );
  NAND2XL U15820 ( .A(n23669), .B(n11403), .Y(n11411) );
  NAND2XL U15821 ( .A(n11402), .B(n11433), .Y(n11403) );
  NOR2XL U15822 ( .A(n11414), .B(n11433), .Y(n11401) );
  NAND2XL U15823 ( .A(n11285), .B(n11284), .Y(n11309) );
  AOI22XL U15824 ( .A0(n7389), .A1(target_temp[27]), .B0(in_valid_d), .B1(
        w1[27]), .Y(n7394) );
  AOI22XL U15825 ( .A0(n6733), .A1(target_temp[28]), .B0(in_valid_d), .B1(
        w1[28]), .Y(n7392) );
  AOI22XL U15826 ( .A0(n7389), .A1(target_temp[29]), .B0(in_valid_d), .B1(
        w1[29]), .Y(n7390) );
  AOI22XL U15827 ( .A0(n6733), .A1(target_temp[26]), .B0(in_valid_d), .B1(
        w1[26]), .Y(n7396) );
  NOR2XL U15828 ( .A(n7847), .B(n7846), .Y(n7851) );
  INVXL U15829 ( .A(n7845), .Y(n7846) );
  INVXL U15830 ( .A(n7848), .Y(n7850) );
  NOR2XL U15831 ( .A(n7841), .B(n7840), .Y(n7844) );
  INVXL U15832 ( .A(n7839), .Y(n7840) );
  NOR2XL U15833 ( .A(n7853), .B(n7852), .Y(n7863) );
  NOR2XL U15834 ( .A(n7859), .B(n7858), .Y(n7860) );
  NOR2XL U15835 ( .A(n7857), .B(n7856), .Y(n7861) );
  NOR2XL U15836 ( .A(n7855), .B(n7854), .Y(n7862) );
  INVXL U15837 ( .A(n10687), .Y(n10688) );
  INVXL U15838 ( .A(n10685), .Y(n10690) );
  INVXL U15839 ( .A(n10684), .Y(n10691) );
  NAND2XL U15840 ( .A(n14427), .B(y10[29]), .Y(n9137) );
  NAND2XL U15841 ( .A(n25233), .B(sigma10[29]), .Y(n9138) );
  NAND2XL U15842 ( .A(n4826), .B(y12[29]), .Y(n9136) );
  INVXL U15843 ( .A(n10677), .Y(n10679) );
  INVXL U15844 ( .A(n10680), .Y(n10682) );
  NAND2XL U15845 ( .A(n9115), .B(n24022), .Y(n9116) );
  NAND2XL U15846 ( .A(n25233), .B(sigma10[23]), .Y(n9115) );
  NAND2XL U15847 ( .A(n14427), .B(y10[25]), .Y(n9123) );
  NAND2XL U15848 ( .A(n25233), .B(sigma10[25]), .Y(n9124) );
  NAND2XL U15849 ( .A(n4826), .B(y12[25]), .Y(n9122) );
  INVXL U15850 ( .A(n10672), .Y(n10673) );
  INVXL U15851 ( .A(n10671), .Y(n10675) );
  AOI22XL U15852 ( .A0(n25233), .A1(data[23]), .B0(in_valid_d), .B1(w1[279]), 
        .Y(n9154) );
  AOI22XL U15853 ( .A0(n25233), .A1(data[24]), .B0(in_valid_d), .B1(w1[280]), 
        .Y(n9152) );
  AOI22XL U15854 ( .A0(n25233), .A1(data[25]), .B0(in_valid_d), .B1(w1[281]), 
        .Y(n9157) );
  AOI22XL U15855 ( .A0(n25233), .A1(data[29]), .B0(in_valid_d), .B1(w1[285]), 
        .Y(n9143) );
  AOI22XL U15856 ( .A0(n4566), .A1(data[30]), .B0(in_valid_d), .B1(w1[286]), 
        .Y(n9140) );
  NAND2XL U15857 ( .A(n3223), .B(learning_rate[30]), .Y(n9141) );
  NAND2XL U15858 ( .A(in_valid_d), .B(w1[155]), .Y(n14438) );
  NAND2XL U15859 ( .A(n25233), .B(learning_rate[27]), .Y(n14439) );
  NAND2XL U15860 ( .A(in_valid_d), .B(w1[156]), .Y(n14434) );
  NAND2XL U15861 ( .A(n25233), .B(learning_rate[28]), .Y(n14435) );
  NAND2XL U15862 ( .A(in_valid_d), .B(w1[158]), .Y(n14403) );
  NAND2XL U15863 ( .A(n25233), .B(learning_rate[30]), .Y(n14404) );
  INVXL U15864 ( .A(n14698), .Y(n14699) );
  INVXL U15865 ( .A(n14697), .Y(n14702) );
  INVXL U15866 ( .A(n14703), .Y(n14708) );
  INVXL U15867 ( .A(n14704), .Y(n14706) );
  NOR2XL U15868 ( .A(n14714), .B(n14713), .Y(n14718) );
  NOR2XL U15869 ( .A(n14712), .B(n14711), .Y(n14719) );
  NOR2XL U15870 ( .A(n14716), .B(n14715), .Y(n14717) );
  NOR2XL U15871 ( .A(n14710), .B(n14709), .Y(n14720) );
  NAND2XL U15872 ( .A(in_valid_t), .B(w2[25]), .Y(n11561) );
  NAND2XL U15873 ( .A(n21166), .B(sigma10[25]), .Y(n11562) );
  NAND2XL U15874 ( .A(n5015), .B(data[57]), .Y(n11563) );
  INVXL U15875 ( .A(n13012), .Y(n13014) );
  NAND2XL U15876 ( .A(in_valid_t), .B(w2[29]), .Y(n11573) );
  NAND2XL U15877 ( .A(n21166), .B(sigma10[29]), .Y(n11574) );
  NAND2XL U15878 ( .A(n5032), .B(data[61]), .Y(n11575) );
  INVXL U15879 ( .A(n13006), .Y(n13008) );
  NOR2XL U15880 ( .A(n13011), .B(n13010), .Y(n13016) );
  INVXL U15881 ( .A(n13009), .Y(n13011) );
  INVXL U15882 ( .A(n17405), .Y(n17407) );
  INVXL U15883 ( .A(n17402), .Y(n17404) );
  INVXL U15884 ( .A(n23498), .Y(n23499) );
  NAND2XL U15885 ( .A(n23915), .B(n23497), .Y(n23500) );
  XOR2XL U15886 ( .A(n23918), .B(n23917), .Y(n23927) );
  INVXL U15887 ( .A(n23916), .Y(n23917) );
  NAND2XL U15888 ( .A(n23915), .B(n23914), .Y(n23918) );
  XOR2XL U15889 ( .A(n23504), .B(n23503), .Y(n23928) );
  NAND2XL U15890 ( .A(n23915), .B(n23502), .Y(n23504) );
  INVXL U15891 ( .A(n23501), .Y(n23502) );
  XOR2XL U15892 ( .A(n23906), .B(n23905), .Y(n23948) );
  NAND2XL U15893 ( .A(n23915), .B(n23904), .Y(n23906) );
  INVXL U15894 ( .A(n23903), .Y(n23904) );
  XOR2XL U15895 ( .A(n20772), .B(n20771), .Y(n23933) );
  NAND2XL U15896 ( .A(n23915), .B(n20770), .Y(n20772) );
  INVXL U15897 ( .A(n20769), .Y(n20770) );
  XOR2XL U15898 ( .A(n23601), .B(n23600), .Y(n23907) );
  INVXL U15899 ( .A(n23599), .Y(n23600) );
  NAND2XL U15900 ( .A(n23915), .B(n23598), .Y(n23601) );
  INVXL U15901 ( .A(n20766), .Y(n20767) );
  NAND2XL U15902 ( .A(n23915), .B(n20765), .Y(n20768) );
  NAND2X1 U15903 ( .A(n3537), .B(n5100), .Y(n23538) );
  XOR2XL U15904 ( .A(n11475), .B(n11474), .Y(n23886) );
  INVXL U15905 ( .A(n11473), .Y(n11474) );
  NAND2XL U15906 ( .A(n23915), .B(n11472), .Y(n11475) );
  XOR2XL U15907 ( .A(n11469), .B(n20293), .Y(n23919) );
  NAND2XL U15908 ( .A(n23915), .B(n11467), .Y(n11469) );
  INVXL U15909 ( .A(n20292), .Y(n11467) );
  XOR2XL U15910 ( .A(n19082), .B(n19081), .Y(n23725) );
  NAND2XL U15911 ( .A(n23915), .B(n19080), .Y(n19082) );
  XOR2XL U15912 ( .A(n23898), .B(n23897), .Y(n23932) );
  INVXL U15913 ( .A(n23896), .Y(n23897) );
  NAND2XL U15914 ( .A(n23915), .B(n23895), .Y(n23898) );
  XOR2XL U15915 ( .A(n23597), .B(n23596), .Y(n23899) );
  NAND2XL U15916 ( .A(n23915), .B(n23595), .Y(n23597) );
  INVXL U15917 ( .A(n23594), .Y(n23595) );
  XOR2XL U15918 ( .A(n11130), .B(n11129), .Y(n20957) );
  NAND2XL U15919 ( .A(n11128), .B(n11127), .Y(n11129) );
  AOI21XL U15920 ( .A0(n11279), .A1(n11277), .B0(n11125), .Y(n11130) );
  INVXL U15921 ( .A(n11126), .Y(n11128) );
  NOR2XL U15922 ( .A(n11461), .B(n11460), .Y(n20958) );
  INVXL U15923 ( .A(n11459), .Y(n11460) );
  NAND2XL U15924 ( .A(n20958), .B(n20957), .Y(n20959) );
  NAND2XL U15925 ( .A(n17367), .B(n17366), .Y(n17368) );
  XNOR2XL U15926 ( .A(n23915), .B(n19063), .Y(n19083) );
  XOR2XL U15927 ( .A(n19067), .B(n20959), .Y(n20962) );
  NAND2XL U15928 ( .A(n19066), .B(n19065), .Y(n19067) );
  INVXL U15929 ( .A(n19064), .Y(n19066) );
  XOR2XL U15930 ( .A(n11379), .B(n11378), .Y(n20721) );
  INVXL U15931 ( .A(n23468), .Y(n23469) );
  NAND2XL U15932 ( .A(n23915), .B(n23467), .Y(n23470) );
  XOR2XL U15933 ( .A(n23466), .B(n23465), .Y(n23885) );
  NAND2XL U15934 ( .A(n23915), .B(n23464), .Y(n23466) );
  INVXL U15935 ( .A(n23463), .Y(n23464) );
  AOI21XL U15936 ( .A0(n18843), .A1(n18842), .B0(n18841), .Y(n18844) );
  XOR2XL U15937 ( .A(n18840), .B(n18839), .Y(n18842) );
  INVXL U15938 ( .A(n20623), .Y(n20294) );
  NAND2XL U15939 ( .A(n23915), .B(n20622), .Y(n20295) );
  INVXL U15940 ( .A(n20625), .Y(n20719) );
  NAND2XL U15941 ( .A(n20623), .B(n20622), .Y(n20718) );
  NOR2XL U15942 ( .A(n20719), .B(n20718), .Y(n20724) );
  XNOR2XL U15943 ( .A(n11095), .B(n11094), .Y(n20725) );
  NAND2XL U15944 ( .A(n11309), .B(n11326), .Y(n11308) );
  NAND2XL U15945 ( .A(n11287), .B(n11286), .Y(n11326) );
  NOR2XL U15946 ( .A(n11404), .B(n23785), .Y(n25713) );
  NOR2XL U15947 ( .A(n11308), .B(n11440), .Y(n11305) );
  NAND2XL U15948 ( .A(n11289), .B(n11288), .Y(n11439) );
  NAND2XL U15949 ( .A(n24443), .B(n24440), .Y(n25831) );
  NAND2XL U15950 ( .A(n25716), .B(n25713), .Y(n25070) );
  NAND2XL U15951 ( .A(n11305), .B(n11439), .Y(n11301) );
  NOR2XL U15952 ( .A(n11405), .B(n25070), .Y(n24440) );
  NOR2XL U15953 ( .A(n11301), .B(n11435), .Y(n11298) );
  NAND2XL U15954 ( .A(n11291), .B(n11290), .Y(n11434) );
  NAND2XL U15955 ( .A(n11298), .B(n11434), .Y(n11294) );
  NAND2BXL U15956 ( .AN(n11402), .B(n11401), .Y(n23669) );
  NOR2XL U15957 ( .A(n11411), .B(n11410), .Y(n23674) );
  NOR2XL U15958 ( .A(n23680), .B(n11409), .Y(n11410) );
  NAND3BXL U15959 ( .AN(n11408), .B(n25835), .C(n24443), .Y(n11409) );
  OR2XL U15960 ( .A(n20570), .B(n20569), .Y(n20571) );
  NAND2XL U15961 ( .A(n24786), .B(n24785), .Y(n24788) );
  INVXL U15962 ( .A(n24784), .Y(n24786) );
  INVXL U15963 ( .A(n25804), .Y(n25806) );
  NAND2XL U15964 ( .A(n20558), .B(n20557), .Y(n20559) );
  INVXL U15965 ( .A(n23616), .Y(n23826) );
  NAND2X1 U15966 ( .A(n20368), .B(n5100), .Y(n5592) );
  INVXL U15967 ( .A(n20369), .Y(n20370) );
  NAND2XL U15968 ( .A(n9172), .B(n9171), .Y(n9173) );
  INVXL U15969 ( .A(n9170), .Y(n9172) );
  INVXL U15970 ( .A(n20801), .Y(n20802) );
  XOR2XL U15971 ( .A(n9178), .B(n9189), .Y(n20791) );
  NAND2XL U15972 ( .A(n9177), .B(n9176), .Y(n9178) );
  INVXL U15973 ( .A(n9175), .Y(n9177) );
  OAI21X2 U15974 ( .A0(n15558), .A1(n14919), .B0(n14918), .Y(n24100) );
  INVXL U15975 ( .A(n24399), .Y(n15741) );
  XOR2XL U15976 ( .A(n9145), .B(n10677), .Y(n9185) );
  INVXL U15977 ( .A(n24384), .Y(n24385) );
  INVXL U15978 ( .A(n24269), .Y(n24267) );
  NOR2XL U15979 ( .A(n20136), .B(n20135), .Y(n24067) );
  INVXL U15980 ( .A(temp1[31]), .Y(n19351) );
  NOR2XL U15981 ( .A(n21111), .B(temp2[31]), .Y(n19348) );
  NAND3XL U15982 ( .A(n3072), .B(n20066), .C(n23200), .Y(n24065) );
  INVXL U15983 ( .A(n20906), .Y(n20903) );
  NOR2XL U15984 ( .A(n20587), .B(n20586), .Y(n20588) );
  INVXL U15985 ( .A(n23805), .Y(n23802) );
  NOR2XL U15986 ( .A(n25352), .B(n23200), .Y(n24570) );
  NAND2X1 U15987 ( .A(n5574), .B(n5100), .Y(n5573) );
  OAI22X1 U15988 ( .A0(n24806), .A1(n24805), .B0(n24804), .B1(n3074), .Y(
        n24860) );
  NOR2XL U15989 ( .A(n24803), .B(n24802), .Y(n24805) );
  NAND2X1 U15990 ( .A(n3132), .B(n20713), .Y(n5526) );
  INVXL U15991 ( .A(n23966), .Y(n23965) );
  NAND3X1 U15992 ( .A(n2988), .B(n23549), .C(n23734), .Y(n5452) );
  NAND2X1 U15993 ( .A(n2988), .B(n23734), .Y(n5450) );
  NAND2XL U15994 ( .A(n3357), .B(n20930), .Y(n20932) );
  NAND2X1 U15995 ( .A(n3357), .B(n5800), .Y(n20746) );
  NOR2X1 U15996 ( .A(n20702), .B(n3015), .Y(n5472) );
  NAND3X1 U15997 ( .A(n4651), .B(n20697), .C(n5771), .Y(n20699) );
  NOR2X1 U15998 ( .A(n14549), .B(n20661), .Y(n14643) );
  NAND2XL U15999 ( .A(n23744), .B(n5388), .Y(n5387) );
  INVXL U16000 ( .A(n20786), .Y(n20658) );
  XOR2XL U16001 ( .A(n14445), .B(n14697), .Y(n14460) );
  XOR2XL U16002 ( .A(n18762), .B(n19032), .Y(n18785) );
  INVXL U16003 ( .A(n6133), .Y(n5912) );
  CMPR32X1 U16004 ( .A(n14715), .B(n24028), .C(n14658), .CO(n24027), .S(n25775) );
  NAND2XL U16005 ( .A(n8482), .B(n8188), .Y(n8162) );
  INVXL U16006 ( .A(n24476), .Y(n24493) );
  NAND2XL U16007 ( .A(n24493), .B(n24492), .Y(n24495) );
  INVXL U16008 ( .A(n24646), .Y(n24627) );
  NOR2XL U16009 ( .A(n24646), .B(n24645), .Y(n24647) );
  INVXL U16010 ( .A(n24725), .Y(n24688) );
  OR2XL U16011 ( .A(n24684), .B(n3075), .Y(n24685) );
  NAND2XL U16012 ( .A(n24754), .B(n24753), .Y(n24755) );
  NAND2XL U16013 ( .A(n24831), .B(n24830), .Y(n24832) );
  NOR2XL U16014 ( .A(n24855), .B(n24854), .Y(n24857) );
  INVXL U16015 ( .A(n24951), .Y(n24903) );
  INVXL U16016 ( .A(n24953), .Y(n24861) );
  NAND2XL U16017 ( .A(n24900), .B(n24899), .Y(n24901) );
  NAND3BXL U16018 ( .AN(n24897), .B(n24896), .C(n3075), .Y(n24900) );
  NAND2BXL U16019 ( .AN(n24996), .B(n24995), .Y(n24997) );
  INVXL U16020 ( .A(n24482), .Y(n24503) );
  INVXL U16021 ( .A(n24518), .Y(n24537) );
  NAND2XL U16022 ( .A(n24585), .B(n24584), .Y(n24587) );
  INVXL U16023 ( .A(n24583), .Y(n24585) );
  INVXL U16024 ( .A(n24637), .Y(n24657) );
  NOR2XL U16025 ( .A(n24658), .B(n24657), .Y(n24659) );
  INVXL U16026 ( .A(n24670), .Y(n24698) );
  NOR2XL U16027 ( .A(n15915), .B(n15914), .Y(n15917) );
  INVXL U16028 ( .A(n24975), .Y(n24928) );
  NAND2X1 U16029 ( .A(in_valid_d), .B(data_point[24]), .Y(n14407) );
  NAND2X1 U16030 ( .A(in_valid_d), .B(data_point[28]), .Y(n14413) );
  NAND2X1 U16031 ( .A(in_valid_d), .B(data_point[30]), .Y(n14416) );
  OAI21X2 U16032 ( .A0(n21628), .A1(n21366), .B0(n21398), .Y(n23402) );
  NAND2XL U16033 ( .A(n23116), .B(n21434), .Y(n21397) );
  NAND2XL U16034 ( .A(n3020), .B(n21413), .Y(n21394) );
  INVXL U16035 ( .A(temp2[31]), .Y(n14966) );
  NOR2XL U16036 ( .A(n21111), .B(temp3[31]), .Y(n14964) );
  NOR2XL U16037 ( .A(n3077), .B(n3076), .Y(n23168) );
  AOI2BB2XL U16038 ( .B0(n22188), .B1(n22222), .A0N(n22222), .A1N(n3126), .Y(
        n23408) );
  INVXL U16039 ( .A(n23409), .Y(n22222) );
  OAI21X2 U16040 ( .A0(n21628), .A1(n21356), .B0(n21399), .Y(n23420) );
  NAND2XL U16041 ( .A(n3020), .B(n21409), .Y(n21395) );
  INVXL U16042 ( .A(n23393), .Y(n22175) );
  NAND3XL U16043 ( .A(n3031), .B(n20597), .C(n8997), .Y(n23175) );
  NOR2XL U16044 ( .A(n21111), .B(temp1[31]), .Y(n8216) );
  NAND2XL U16045 ( .A(n5480), .B(target_temp[25]), .Y(n11594) );
  NAND2XL U16046 ( .A(n5032), .B(sigma10[25]), .Y(n11595) );
  NAND2XL U16047 ( .A(in_valid_t), .B(w2[89]), .Y(n17163) );
  NAND2XL U16048 ( .A(n3111), .B(data[121]), .Y(n17165) );
  NAND2XL U16049 ( .A(n21166), .B(target_temp[28]), .Y(n11582) );
  NAND2XL U16050 ( .A(n5032), .B(sigma10[28]), .Y(n11583) );
  NAND2XL U16051 ( .A(n21166), .B(target_temp[29]), .Y(n11578) );
  NAND2XL U16052 ( .A(n5015), .B(sigma10[29]), .Y(n11579) );
  NAND2XL U16053 ( .A(in_valid_t), .B(w2[93]), .Y(n17176) );
  NAND2XL U16054 ( .A(n4875), .B(data[125]), .Y(n17178) );
  NOR2BX1 U16055 ( .AN(n23638), .B(n23637), .Y(n23640) );
  NAND4XL U16056 ( .A(n19040), .B(n19039), .C(n19038), .D(n19037), .Y(n19041)
         );
  NOR2XL U16057 ( .A(n19036), .B(n19035), .Y(n19037) );
  NAND3XL U16058 ( .A(n22480), .B(n22479), .C(n22478), .Y(n22483) );
  NAND2XL U16059 ( .A(in_valid_t), .B(w2[63]), .Y(n22478) );
  INVXL U16060 ( .A(n25701), .Y(n23716) );
  NAND2XL U16061 ( .A(n23715), .B(n23716), .Y(n23784) );
  NAND2XL U16062 ( .A(n25829), .B(n23675), .Y(n23676) );
  NOR2BXL U16063 ( .AN(n23674), .B(n23673), .Y(n23675) );
  NOR2XL U16064 ( .A(n25832), .B(n25704), .Y(n25700) );
  AOI21XL U16065 ( .A0(n11440), .A1(n11308), .B0(n11305), .Y(n11323) );
  XOR2XL U16066 ( .A(n7399), .B(n7839), .Y(n7411) );
  NAND2XL U16067 ( .A(n9160), .B(n9179), .Y(n9180) );
  NOR2X1 U16068 ( .A(n11412), .B(n11411), .Y(n23668) );
  NOR2XL U16069 ( .A(n11406), .B(n25831), .Y(n23677) );
  INVXL U16070 ( .A(n25832), .Y(n23715) );
  INVXL U16071 ( .A(n7869), .Y(n7388) );
  NAND2XL U16072 ( .A(n11315), .B(n11314), .Y(n11433) );
  NAND2XL U16073 ( .A(n11304), .B(n11303), .Y(n11426) );
  NAND2XL U16074 ( .A(n11300), .B(n11299), .Y(n11427) );
  NAND2XL U16075 ( .A(n11297), .B(n11296), .Y(n11420) );
  NAND2XL U16076 ( .A(n11293), .B(n11292), .Y(n11421) );
  NAND2XL U16077 ( .A(n11283), .B(n11282), .Y(n11418) );
  NAND2XL U16078 ( .A(n11281), .B(n11280), .Y(n11419) );
  MXI2XL U16079 ( .A(n23193), .B(data_point[31]), .S0(n3123), .Y(n23194) );
  NOR4BXL U16080 ( .AN(n10676), .B(n10675), .C(n10674), .D(n10673), .Y(n10702)
         );
  NOR3XL U16081 ( .A(n10683), .B(n10682), .C(n10681), .Y(n10701) );
  NAND4XL U16082 ( .A(n10691), .B(n10690), .C(n10689), .D(n10688), .Y(n10700)
         );
  NAND4XL U16083 ( .A(n10684), .B(n10685), .C(n10686), .D(n10687), .Y(n10668)
         );
  NAND4XL U16084 ( .A(n10694), .B(n10695), .C(n10693), .D(n10692), .Y(n10667)
         );
  NAND2XL U16085 ( .A(in_valid_d), .B(w1[287]), .Y(n25234) );
  NAND2XL U16086 ( .A(n4856), .B(y12[31]), .Y(n25231) );
  NAND2XL U16087 ( .A(n25233), .B(sigma10[31]), .Y(n25232) );
  NAND2XL U16088 ( .A(in_valid_d), .B(data_point[31]), .Y(n25230) );
  NAND4XL U16089 ( .A(n14720), .B(n14719), .C(n14718), .D(n14717), .Y(n14721)
         );
  NAND4XL U16090 ( .A(n14708), .B(n14707), .C(n14706), .D(n14705), .Y(n14722)
         );
  NAND4XL U16091 ( .A(n14702), .B(n14701), .C(n14700), .D(n14699), .Y(n14723)
         );
  NAND2XL U16092 ( .A(n4826), .B(target_temp[31]), .Y(n25236) );
  NAND4XL U16093 ( .A(n13018), .B(n13017), .C(n13016), .D(n13015), .Y(n13023)
         );
  NOR2XL U16094 ( .A(n13008), .B(n13007), .Y(n13017) );
  NOR2XL U16095 ( .A(n13014), .B(n13013), .Y(n13015) );
  INVXL U16096 ( .A(n22484), .Y(n23084) );
  INVXL U16097 ( .A(learning_rate[3]), .Y(n23999) );
  INVXL U16098 ( .A(learning_rate[10]), .Y(n23992) );
  OAI22XL U16099 ( .A0(n25813), .A1(n26310), .B0(n4860), .B1(n25992), .Y(
        n22484) );
  INVX1 U16100 ( .A(n20315), .Y(n20316) );
  NAND2X1 U16101 ( .A(n3895), .B(n20317), .Y(n4928) );
  NOR2XL U16102 ( .A(n23545), .B(n3115), .Y(n23546) );
  NAND2XL U16103 ( .A(n25723), .B(temp0[17]), .Y(n4820) );
  NOR2XL U16104 ( .A(n23941), .B(n9146), .Y(n23942) );
  NOR2XL U16105 ( .A(n11476), .B(n9146), .Y(n11477) );
  CLKINVX3 U16106 ( .A(n2982), .Y(n23884) );
  NAND2X1 U16107 ( .A(n3353), .B(n25298), .Y(n4954) );
  NOR2XL U16108 ( .A(in_valid_d), .B(n25886), .Y(n10719) );
  NOR2XL U16109 ( .A(n23471), .B(n3115), .Y(n23473) );
  NAND2XL U16110 ( .A(n25723), .B(temp0[20]), .Y(n20629) );
  XOR2XL U16111 ( .A(n20626), .B(n20719), .Y(n25725) );
  NAND2XL U16112 ( .A(n23915), .B(n20624), .Y(n20626) );
  INVXL U16113 ( .A(n20718), .Y(n20624) );
  NAND2X1 U16114 ( .A(n3357), .B(n5717), .Y(n20342) );
  INVXL U16115 ( .A(n11302), .Y(n11321) );
  AOI21XL U16116 ( .A0(n11437), .A1(n11294), .B0(n11414), .Y(n11317) );
  AOI21XL U16117 ( .A0(n11435), .A1(n11301), .B0(n11298), .Y(n11329) );
  INVXL U16118 ( .A(n11295), .Y(n11319) );
  AOI22XL U16119 ( .A0(n20385), .A1(n25301), .B0(n25300), .B1(n25299), .Y(
        n25689) );
  INVXL U16120 ( .A(n25301), .Y(n25299) );
  AOI22X1 U16121 ( .A0(n20385), .A1(n23583), .B0(n25300), .B1(n23582), .Y(
        n23768) );
  NOR2XL U16122 ( .A(n3024), .B(n23973), .Y(n25741) );
  OAI2BB1X2 U16123 ( .A0N(n24174), .A1N(n3353), .B0(n4977), .Y(n4976) );
  NAND2X1 U16124 ( .A(n3131), .B(n24183), .Y(n4977) );
  AOI22X1 U16125 ( .A0(n20385), .A1(n20635), .B0(n25300), .B1(n20634), .Y(
        n23841) );
  AOI22X1 U16126 ( .A0(n20385), .A1(n20608), .B0(n25300), .B1(n20607), .Y(
        n25826) );
  INVXL U16127 ( .A(n20608), .Y(n20605) );
  AOI22X1 U16128 ( .A0(n20385), .A1(n20841), .B0(n25300), .B1(n20840), .Y(
        n24675) );
  INVXL U16129 ( .A(n24389), .Y(n24393) );
  INVXL U16130 ( .A(n24432), .Y(n24438) );
  INVXL U16131 ( .A(n24299), .Y(n24303) );
  INVX1 U16132 ( .A(data_point[21]), .Y(n5008) );
  NOR2X1 U16133 ( .A(n4582), .B(n6235), .Y(n25141) );
  INVX1 U16134 ( .A(data_point[13]), .Y(n6285) );
  NOR2X2 U16135 ( .A(n4583), .B(n6154), .Y(n25155) );
  INVX1 U16136 ( .A(data_point[17]), .Y(n6154) );
  INVX1 U16137 ( .A(data_point[22]), .Y(n6271) );
  NOR2X1 U16138 ( .A(n6250), .B(n4584), .Y(n25150) );
  INVX1 U16139 ( .A(data_point[14]), .Y(n6258) );
  INVX1 U16140 ( .A(data_point[16]), .Y(n6267) );
  AOI22X1 U16141 ( .A0(n20385), .A1(n20889), .B0(n25300), .B1(n20888), .Y(
        n23699) );
  INVXL U16142 ( .A(n24340), .Y(n24344) );
  INVXL U16143 ( .A(n24308), .Y(n24312) );
  INVXL U16144 ( .A(n24068), .Y(n24075) );
  INVX1 U16145 ( .A(n20997), .Y(n25577) );
  AOI22XL U16146 ( .A0(n24692), .A1(n20996), .B0(n24908), .B1(n20995), .Y(
        n20997) );
  XOR2XL U16147 ( .A(n24572), .B(n24527), .Y(n20995) );
  AOI22XL U16148 ( .A0(n24692), .A1(n24531), .B0(n24908), .B1(n24530), .Y(
        n24532) );
  INVX1 U16149 ( .A(n24578), .Y(n25545) );
  INVXL U16150 ( .A(n24577), .Y(n24574) );
  AOI22XL U16151 ( .A0(n22486), .A1(sigma11[7]), .B0(n25754), .B1(sigma12[7]), 
        .Y(n24150) );
  NAND2X1 U16152 ( .A(n3895), .B(n21023), .Y(n4931) );
  AOI22X1 U16153 ( .A0(n25503), .A1(n4215), .B0(n4220), .B1(n25527), .Y(n24157) );
  AOI22X1 U16154 ( .A0(n5336), .A1(n20747), .B0(n21052), .B1(n3136), .Y(n24122) );
  AOI22X1 U16155 ( .A0(n20935), .A1(n3136), .B0(n5336), .B1(n20936), .Y(n23697) );
  NOR2XL U16156 ( .A(n20373), .B(cs[2]), .Y(n17459) );
  INVXL U16157 ( .A(n23857), .Y(n23861) );
  INVXL U16158 ( .A(n24294), .Y(n24298) );
  INVXL U16159 ( .A(n23759), .Y(n23763) );
  INVXL U16160 ( .A(n24607), .Y(n24596) );
  INVX1 U16161 ( .A(n24498), .Y(n25596) );
  AOI22XL U16162 ( .A0(n24692), .A1(n24497), .B0(n24908), .B1(n24496), .Y(
        n24498) );
  INVXL U16163 ( .A(n24497), .Y(n24494) );
  AOI22XL U16164 ( .A0(n24692), .A1(n24651), .B0(n24908), .B1(n24650), .Y(
        n24652) );
  INVXL U16165 ( .A(n24651), .Y(n24648) );
  INVX1 U16166 ( .A(n25363), .Y(n25821) );
  AOI22XL U16167 ( .A0(n24692), .A1(n25362), .B0(n24908), .B1(n25361), .Y(
        n25363) );
  INVXL U16168 ( .A(n25362), .Y(n25359) );
  INVXL U16169 ( .A(n14407), .Y(n25218) );
  INVXL U16170 ( .A(n14410), .Y(n25215) );
  INVXL U16171 ( .A(n14413), .Y(n25212) );
  INVXL U16172 ( .A(n14416), .Y(n24021) );
  INVXL U16173 ( .A(n23275), .Y(n23273) );
  XNOR2XL U16174 ( .A(n23288), .B(n23287), .Y(n23289) );
  INVXL U16175 ( .A(n23290), .Y(n23288) );
  INVXL U16176 ( .A(n23242), .Y(n23239) );
  AND3XL U16177 ( .A(n23132), .B(n23131), .C(n23130), .Y(n23137) );
  INVXL U16178 ( .A(n23225), .Y(n23132) );
  INVXL U16179 ( .A(n23282), .Y(n23279) );
  XOR2XL U16180 ( .A(n23293), .B(n23292), .Y(n23284) );
  INVXL U16181 ( .A(n23297), .Y(n23294) );
  INVXL U16182 ( .A(n23265), .Y(n23262) );
  INVXL U16183 ( .A(n23318), .Y(n23245) );
  INVXL U16184 ( .A(n23322), .Y(n23319) );
  NAND2XL U16185 ( .A(n23346), .B(n23313), .Y(n23314) );
  INVXL U16186 ( .A(n23350), .Y(n23347) );
  NAND2XL U16187 ( .A(n23346), .B(n23337), .Y(n23339) );
  INVXL U16188 ( .A(n23311), .Y(n23308) );
  INVXL U16189 ( .A(n23335), .Y(n23332) );
  INVXL U16190 ( .A(n23305), .Y(n23302) );
  INVXL U16191 ( .A(n23376), .Y(n23326) );
  INVXL U16192 ( .A(n23380), .Y(n23377) );
  NAND2XL U16193 ( .A(n23383), .B(n23370), .Y(n23372) );
  INVXL U16194 ( .A(n23387), .Y(n23384) );
  AOI22XL U16195 ( .A0(n23419), .A1(n23230), .B0(n23418), .B1(n23229), .Y(
        n23231) );
  INVXL U16196 ( .A(n23415), .Y(n23233) );
  INVXL U16197 ( .A(learning_rate[8]), .Y(n23994) );
  INVXL U16198 ( .A(learning_rate[17]), .Y(n23989) );
  INVXL U16199 ( .A(learning_rate[24]), .Y(n23980) );
  INVXL U16200 ( .A(learning_rate[25]), .Y(n24006) );
  INVXL U16201 ( .A(learning_rate[27]), .Y(n23053) );
  NAND2XL U16202 ( .A(n24015), .B(n24011), .Y(n24007) );
  NAND2BXL U16203 ( .AN(n23976), .B(n24012), .Y(n24008) );
  OAI22XL U16204 ( .A0(n22482), .A1(n22481), .B0(n22483), .B1(n22484), .Y(
        n25258) );
  NOR2XL U16205 ( .A(n22485), .B(n23084), .Y(n25257) );
  INVXL U16206 ( .A(n22483), .Y(n22485) );
  OAI211XL U16207 ( .A0(n23716), .A1(n25829), .B0(n23784), .C0(n25699), .Y(
        n23717) );
  AOI21XL U16208 ( .A0(n23868), .A1(n23718), .B0(n23863), .Y(n5357) );
  NAND2X1 U16209 ( .A(n23864), .B(n23862), .Y(n5358) );
  INVXL U16210 ( .A(n23678), .Y(n23680) );
  INVXL U16211 ( .A(temp0[31]), .Y(n25246) );
  INVX1 U16212 ( .A(n25723), .Y(n25837) );
  OAI22XL U16213 ( .A0(n11446), .A1(n11445), .B0(n11444), .B1(n11443), .Y(
        n25244) );
  AOI21XL U16214 ( .A0(n23199), .A1(n23198), .B0(n23197), .Y(n25691) );
  XOR2XL U16215 ( .A(n23196), .B(n23195), .Y(n23197) );
  AOI22XL U16216 ( .A0(n6733), .A1(target_temp[31]), .B0(in_valid_d), .B1(
        w1[31]), .Y(n23196) );
  OAI21XL U16217 ( .A0(n25241), .A1(n25240), .B0(n25239), .Y(n25660) );
  XOR2XL U16218 ( .A(n25238), .B(n25237), .Y(n25239) );
  NAND3XL U16219 ( .A(n25232), .B(n25231), .C(n25230), .Y(n25238) );
  NAND3XL U16220 ( .A(n25236), .B(n25235), .C(n25234), .Y(n25237) );
  NOR2XL U16221 ( .A(n23084), .B(n23083), .Y(n25666) );
  OAI2BB1XL U16222 ( .A0N(n22477), .A1N(n24036), .B0(n22476), .Y(n25670) );
  XNOR2XL U16223 ( .A(n22475), .B(n22474), .Y(n22476) );
  AOI22XL U16224 ( .A0(n23082), .A1(n23081), .B0(n23083), .B1(n23084), .Y(
        n25668) );
  INVXL U16225 ( .A(n23078), .Y(n23081) );
  INVXL U16226 ( .A(n24050), .Y(n23082) );
  INVXL U16227 ( .A(n23970), .Y(n23049) );
  NOR3XL U16228 ( .A(n25541), .B(n23072), .C(n23071), .Y(n2489) );
  NAND2X1 U16229 ( .A(n17430), .B(n5336), .Y(n5833) );
  NAND2X1 U16230 ( .A(n17439), .B(n3136), .Y(n5832) );
  OAI21XL U16231 ( .A0(n25093), .A1(n4581), .B0(n24278), .Y(n2563) );
  OAI21XL U16232 ( .A0(n24449), .A1(n4581), .B0(n24398), .Y(n2561) );
  OAI2BB1XL U16233 ( .A0N(n25807), .A1N(n20785), .B0(n20784), .Y(n2565) );
  AOI2BB2X1 U16234 ( .B0(n2983), .B1(temp2[26]), .A0N(n25722), .A1N(n4582), 
        .Y(n20784) );
  NAND2XL U16235 ( .A(n25723), .B(temp0[7]), .Y(n23921) );
  OAI21XL U16236 ( .A0(n24616), .A1(n3121), .B0(n23510), .Y(n2598) );
  NAND2XL U16237 ( .A(n25723), .B(temp0[9]), .Y(n23506) );
  AOI21XL U16238 ( .A0(n24644), .A1(in_valid_d), .B0(n23953), .Y(n23954) );
  NAND2BXL U16239 ( .AN(n23952), .B(n23951), .Y(n23953) );
  NAND2XL U16240 ( .A(n25723), .B(temp0[10]), .Y(n23951) );
  OAI21XL U16241 ( .A0(n3121), .A1(n20844), .B0(n6005), .Y(n2533) );
  INVXL U16242 ( .A(n17440), .Y(mul5_out[10]) );
  NAND2X1 U16243 ( .A(n17430), .B(n3136), .Y(n5707) );
  OAI211XL U16244 ( .A0(n24868), .A1(n4582), .B0(n19046), .C0(n19045), .Y(
        n2581) );
  OAI211XL U16245 ( .A0(n24735), .A1(n4586), .B0(n19052), .C0(n19051), .Y(
        n2589) );
  NAND2XL U16246 ( .A(n25723), .B(temp0[8]), .Y(n4844) );
  NAND2BXL U16247 ( .AN(n23729), .B(n23728), .Y(n23730) );
  NAND2XL U16248 ( .A(n25723), .B(temp0[3]), .Y(n23728) );
  NAND2XL U16249 ( .A(n25723), .B(temp0[14]), .Y(n23935) );
  NAND2XL U16250 ( .A(n25723), .B(temp0[11]), .Y(n23909) );
  OAI2BB1XL U16251 ( .A0N(n25807), .A1N(n20776), .B0(n20775), .Y(n2586) );
  NAND2XL U16252 ( .A(n25723), .B(temp0[15]), .Y(n4824) );
  NAND3XL U16253 ( .A(n2990), .B(n23654), .C(n23653), .Y(n2541) );
  NAND3BXL U16254 ( .AN(n4836), .B(n23705), .C(n23704), .Y(n2538) );
  NOR2XL U16255 ( .A(n23602), .B(n3115), .Y(n23603) );
  NAND2XL U16256 ( .A(n25723), .B(temp0[5]), .Y(n23888) );
  OAI21XL U16257 ( .A0(n24821), .A1(n3121), .B0(n20827), .Y(n2584) );
  NAND2XL U16258 ( .A(n25723), .B(temp0[16]), .Y(n4873) );
  NAND2XL U16259 ( .A(n25723), .B(temp0[6]), .Y(n5103) );
  OR2X2 U16260 ( .A(n24190), .B(n3121), .Y(n5207) );
  NAND2X1 U16261 ( .A(n23795), .B(n5366), .Y(n20978) );
  OAI2BB1XL U16262 ( .A0N(n19089), .A1N(n25807), .B0(n19088), .Y(n2612) );
  NAND2BXL U16263 ( .AN(n19086), .B(n19085), .Y(n19087) );
  NAND2XL U16264 ( .A(n25723), .B(temp0[2]), .Y(n19085) );
  NAND2XL U16265 ( .A(n25723), .B(temp0[13]), .Y(n4846) );
  NAND2XL U16266 ( .A(n25723), .B(temp0[0]), .Y(n4841) );
  NAND2X1 U16267 ( .A(n3001), .B(n3136), .Y(n4866) );
  AOI211X1 U16268 ( .A0(n25723), .A1(temp0[1]), .B0(n19070), .C0(n19069), .Y(
        n19071) );
  NOR2XL U16269 ( .A(n19068), .B(n3115), .Y(n19069) );
  NOR2XL U16270 ( .A(n23770), .B(n4582), .Y(n19070) );
  NOR2XL U16271 ( .A(n23884), .B(n26564), .Y(n4716) );
  AOI21X1 U16272 ( .A0(n25828), .A1(in_valid_d), .B0(n20731), .Y(n20732) );
  OAI2BB1XL U16273 ( .A0N(n25728), .A1N(n20730), .B0(n20729), .Y(n20731) );
  INVX1 U16274 ( .A(n19089), .Y(n24481) );
  NAND2XL U16275 ( .A(n5967), .B(n25807), .Y(n5951) );
  OAI211XL U16276 ( .A0(n24224), .A1(n4585), .B0(n20675), .C0(n20674), .Y(
        n2537) );
  OAI211XL U16277 ( .A0(n24744), .A1(n4583), .B0(n20314), .C0(n20313), .Y(
        n2539) );
  OAI21XL U16278 ( .A0(n24053), .A1(n4584), .B0(n24052), .Y(n2525) );
  OAI21XL U16279 ( .A0(n25681), .A1(n4586), .B0(n25680), .Y(n2528) );
  OAI21XL U16280 ( .A0(n24290), .A1(n4582), .B0(n24289), .Y(n2527) );
  OAI21XL U16281 ( .A0(n25799), .A1(n4585), .B0(n25798), .Y(n2524) );
  OAI21XL U16282 ( .A0(n25809), .A1(n4583), .B0(n25808), .Y(n2531) );
  AOI22XL U16283 ( .A0(n25378), .A1(n25636), .B0(temp2[19]), .B1(n2984), .Y(
        n23567) );
  NAND2BX1 U16284 ( .AN(n20630), .B(n20629), .Y(n20631) );
  NAND2X1 U16285 ( .A(n5336), .B(n20935), .Y(n6044) );
  OAI21XL U16286 ( .A0(n25709), .A1(n3121), .B0(n25708), .Y(n2568) );
  OAI22XL U16287 ( .A0(n25705), .A1(n3115), .B0(n25837), .B1(n26545), .Y(
        n25706) );
  OAI21XL U16288 ( .A0(n25722), .A1(n3121), .B0(n25721), .Y(n2564) );
  OAI22XL U16289 ( .A0(n25718), .A1(n3115), .B0(n25837), .B1(n26546), .Y(
        n25719) );
  AOI211XL U16290 ( .A0(n25717), .A1(n25716), .B0(n25834), .C0(n25715), .Y(
        n25718) );
  OAI21XL U16291 ( .A0(n25842), .A1(n3121), .B0(n25841), .Y(n2558) );
  OAI22XL U16292 ( .A0(n25838), .A1(n3115), .B0(n25837), .B1(n26594), .Y(
        n25839) );
  AOI211XL U16293 ( .A0(n25836), .A1(n25835), .B0(n25834), .C0(n25833), .Y(
        n25838) );
  OAI21XL U16294 ( .A0(n25093), .A1(n3121), .B0(n25077), .Y(n2562) );
  OAI22XL U16295 ( .A0(n25074), .A1(n3115), .B0(n25837), .B1(n26515), .Y(
        n25075) );
  AOI211XL U16296 ( .A0(n25073), .A1(n25072), .B0(n25834), .C0(n25071), .Y(
        n25074) );
  OAI21XL U16297 ( .A0(n24449), .A1(n3121), .B0(n24448), .Y(n2560) );
  OAI22XL U16298 ( .A0(n24445), .A1(n3115), .B0(n25837), .B1(n26514), .Y(
        n24446) );
  AOI211XL U16299 ( .A0(n24444), .A1(n24443), .B0(n25834), .C0(n24442), .Y(
        n24445) );
  OAI21XL U16300 ( .A0(n9039), .A1(n3227), .B0(n9038), .Y(n9040) );
  AOI22XL U16301 ( .A0(n25025), .A1(y10[28]), .B0(n3050), .B1(y12[28]), .Y(
        n9038) );
  AOI22XL U16302 ( .A0(n25025), .A1(y10[17]), .B0(n8104), .B1(y12[17]), .Y(
        n23609) );
  AOI22XL U16303 ( .A0(n24739), .A1(y12[12]), .B0(n3050), .B1(y11[12]), .Y(
        n24671) );
  AOI22XL U16304 ( .A0(n25025), .A1(y10[15]), .B0(n25656), .B1(y12[15]), .Y(
        n24794) );
  AOI22XL U16305 ( .A0(n22486), .A1(sigma11[27]), .B0(sigma12[27]), .B1(n25754), .Y(n25172) );
  OAI21XL U16306 ( .A0(n25709), .A1(n24632), .B0(n24096), .Y(n24097) );
  AOI22XL U16307 ( .A0(n25025), .A1(y12[19]), .B0(n3050), .B1(y11[19]), .Y(
        n24933) );
  AOI22XL U16308 ( .A0(n25815), .A1(y10[5]), .B0(n25656), .B1(y12[5]), .Y(
        n24545) );
  AOI22XL U16309 ( .A0(n25815), .A1(y10[2]), .B0(n3050), .B1(y12[2]), .Y(
        n24487) );
  AOI22XL U16310 ( .A0(n25815), .A1(y10[1]), .B0(n25656), .B1(y12[1]), .Y(
        n24472) );
  AOI22XL U16311 ( .A0(n25815), .A1(y12[6]), .B0(n25656), .B1(y11[6]), .Y(
        n24559) );
  AOI22XL U16312 ( .A0(n25025), .A1(y12[29]), .B0(n3120), .B1(y11[29]), .Y(
        n25102) );
  AOI22XL U16313 ( .A0(n25815), .A1(y10[25]), .B0(n3050), .B1(y12[25]), .Y(
        n24422) );
  AOI22XL U16314 ( .A0(n25025), .A1(y10[24]), .B0(n3050), .B1(y12[24]), .Y(
        n23876) );
  AOI22XL U16315 ( .A0(n25815), .A1(y12[27]), .B0(n3120), .B1(y11[27]), .Y(
        n25094) );
  AOI21XL U16316 ( .A0(n25220), .A1(n23646), .B0(n25219), .Y(n23647) );
  OAI21XL U16317 ( .A0(n25435), .A1(n4574), .B0(n25434), .Y(n2073) );
  AOI22XL U16318 ( .A0(n3052), .A1(n26135), .B0(n3061), .B1(n26468), .Y(n25434) );
  AOI21XL U16319 ( .A0(n23044), .A1(n23043), .B0(n23042), .Y(n2254) );
  OAI2BB1XL U16320 ( .A0N(n23041), .A1N(n23043), .B0(n23040), .Y(n23042) );
  AOI22XL U16321 ( .A0(n23428), .A1(target_temp[22]), .B0(in_valid_t), .B1(
        target[22]), .Y(n23040) );
  INVXL U16322 ( .A(n25691), .Y(n25694) );
  AOI22XL U16323 ( .A0(n4575), .A1(n26318), .B0(n3061), .B1(n26049), .Y(n25251) );
  AOI22XL U16324 ( .A0(n25820), .A1(n26048), .B0(in_valid_w2), .B1(n26314), 
        .Y(n25682) );
  OAI2BB1XL U16325 ( .A0N(w1[383]), .A1N(n25410), .B0(n25252), .Y(n25253) );
  AOI22XL U16326 ( .A0(n3028), .A1(w1[287]), .B0(in_valid_w1), .B1(weight1[31]), .Y(n25252) );
  AOI22XL U16327 ( .A0(n25815), .A1(y12[31]), .B0(n25656), .B1(y11[31]), .Y(
        n25657) );
  AOI22XL U16328 ( .A0(n25661), .A1(n3050), .B0(y11[31]), .B1(n24958), .Y(
        n25662) );
  INVXL U16329 ( .A(n25660), .Y(n25661) );
  AOI222XL U16330 ( .A0(n25665), .A1(n25292), .B0(w2[63]), .B1(n25820), .C0(
        w2[95]), .C1(in_valid_w2), .Y(n2199) );
  AOI22XL U16331 ( .A0(n4575), .A1(n26049), .B0(n3061), .B1(n26377), .Y(n25250) );
  AOI31XL U16332 ( .A0(n25668), .A1(n25767), .A2(n23087), .B0(n23086), .Y(
        n2295) );
  INVXL U16333 ( .A(n25666), .Y(n23087) );
  AOI22XL U16334 ( .A0(n22486), .A1(sigma11[31]), .B0(n25754), .B1(sigma12[31]), .Y(n23085) );
  AOI21XL U16335 ( .A0(n25754), .A1(n22489), .B0(n22488), .Y(n2359) );
  OAI31XL U16336 ( .A0(n25258), .A1(n3111), .A2(n25257), .B0(n22487), .Y(
        n22488) );
  INVXL U16337 ( .A(n25670), .Y(n22489) );
  AOI22XL U16338 ( .A0(n22486), .A1(sigma12[31]), .B0(n25750), .B1(sigma11[31]), .Y(n22487) );
  MXI2XL U16339 ( .A(mul5_out[31]), .B(n25256), .S0(n5015), .Y(n2358) );
  OAI22XL U16340 ( .A0(n25255), .A1(n26067), .B0(n3050), .B1(n26316), .Y(
        n25256) );
  AOI222XL U16341 ( .A0(n23088), .A1(w1[81]), .B0(n21113), .B1(w1[49]), .C0(
        w1[177]), .C1(n3216), .Y(n1820) );
  AOI222XL U16342 ( .A0(n23088), .A1(w1[211]), .B0(n4577), .B1(w1[179]), .C0(
        w1[307]), .C1(n3216), .Y(n1956) );
  AOI222XL U16343 ( .A0(n3061), .A1(w1[208]), .B0(n4578), .B1(w1[176]), .C0(
        w1[304]), .C1(n3216), .Y(n1944) );
  AOI222XL U16344 ( .A0(n3061), .A1(w1[112]), .B0(n4578), .B1(w1[80]), .C0(
        w1[208]), .C1(n3216), .Y(n1817) );
  AOI22XL U16345 ( .A0(n4575), .A1(n26073), .B0(n23088), .B1(n26366), .Y(
        n25575) );
  AOI22XL U16346 ( .A0(n3052), .A1(n26039), .B0(n3061), .B1(n26367), .Y(n25605) );
  AOI22XL U16347 ( .A0(n3052), .A1(n26097), .B0(n23088), .B1(n26407), .Y(
        n25587) );
  AOI22XL U16348 ( .A0(n3052), .A1(n26027), .B0(n3061), .B1(n26368), .Y(n25619) );
  AOI22XL U16349 ( .A0(n3052), .A1(n26321), .B0(n23088), .B1(n26052), .Y(
        n25616) );
  AOI22XL U16350 ( .A0(n3052), .A1(n26053), .B0(n25542), .B1(n26400), .Y(
        n25650) );
  AOI22XL U16351 ( .A0(n4575), .A1(n26081), .B0(n25542), .B1(n26399), .Y(
        n25629) );
  AOI22XL U16352 ( .A0(n3023), .A1(n26315), .B0(n3061), .B1(n26058), .Y(n25493) );
  AOI22XL U16353 ( .A0(n3052), .A1(n26320), .B0(n3061), .B1(n26051), .Y(n25478) );
  AOI22XL U16354 ( .A0(n25410), .A1(n26058), .B0(n3061), .B1(n26362), .Y(
        n25492) );
  AOI22XL U16355 ( .A0(n4575), .A1(n26080), .B0(n3061), .B1(n26396), .Y(n25583) );
  AOI22XL U16356 ( .A0(n4575), .A1(n26070), .B0(n26353), .B1(n3061), .Y(n25117) );
  AOI22XL U16357 ( .A0(n4575), .A1(n26324), .B0(n3061), .B1(n26057), .Y(n25228) );
  AOI22XL U16358 ( .A0(n4575), .A1(n26078), .B0(n3061), .B1(n26394), .Y(n25563) );
  AOI22XL U16359 ( .A0(n4575), .A1(n26091), .B0(n3061), .B1(n26393), .Y(n25551) );
  AOI22XL U16360 ( .A0(n4575), .A1(n26102), .B0(n3061), .B1(n26376), .Y(n25225) );
  AOI22XL U16361 ( .A0(n3052), .A1(n26072), .B0(n3061), .B1(n26365), .Y(n25468) );
  AOI22XL U16362 ( .A0(n3023), .A1(n26088), .B0(n3061), .B1(n26390), .Y(n25514) );
  AOI22XL U16363 ( .A0(n25410), .A1(n26087), .B0(n3061), .B1(n26389), .Y(
        n25501) );
  AOI22XL U16364 ( .A0(n3052), .A1(n26085), .B0(n23088), .B1(n26385), .Y(
        n25453) );
  AOI22XL U16365 ( .A0(n3023), .A1(n26103), .B0(n3061), .B1(n26378), .Y(n25254) );
  AOI22XL U16366 ( .A0(n4575), .A1(n26105), .B0(n3061), .B1(n26363), .Y(n25516) );
  AOI22XL U16367 ( .A0(n3023), .A1(n26052), .B0(n3061), .B1(n26398), .Y(n25615) );
  AOI22XL U16368 ( .A0(n4575), .A1(n26092), .B0(n23088), .B1(n26397), .Y(
        n25602) );
  INVXL U16369 ( .A(n21171), .Y(n21172) );
  AOI222XL U16370 ( .A0(n3216), .A1(w1[380]), .B0(n21113), .B1(w1[252]), .C0(
        w1[284]), .C1(in_valid_w1), .Y(n21171) );
  AOI22XL U16371 ( .A0(n3023), .A1(n26095), .B0(n3061), .B1(n26405), .Y(n25564) );
  AOI22XL U16372 ( .A0(n3052), .A1(n26068), .B0(n3061), .B1(n26354), .Y(n25653) );
  AOI22XL U16373 ( .A0(n3052), .A1(n26059), .B0(n3061), .B1(n26401), .Y(n25698) );
  AOI22XL U16374 ( .A0(n3052), .A1(n26051), .B0(n25542), .B1(n26387), .Y(
        n25477) );
  AOI22XL U16375 ( .A0(n3052), .A1(n26086), .B0(n3061), .B1(n26386), .Y(n25465) );
  AOI22XL U16376 ( .A0(n3023), .A1(n26075), .B0(n3061), .B1(n26409), .Y(n25652) );
  AOI22XL U16377 ( .A0(n3028), .A1(w1[3]), .B0(in_valid_w1), .B1(w1[131]), .Y(
        n25606) );
  AOI22XL U16378 ( .A0(n3028), .A1(w1[2]), .B0(in_valid_w1), .B1(w1[130]), .Y(
        n25620) );
  AOI22XL U16379 ( .A0(n3064), .A1(w1[8]), .B0(in_valid_w1), .B1(w1[136]), .Y(
        n21126) );
  AOI22XL U16380 ( .A0(n3028), .A1(w1[11]), .B0(in_valid_w1), .B1(w1[139]), 
        .Y(n21132) );
  AOI22XL U16381 ( .A0(n3064), .A1(w1[12]), .B0(in_valid_w1), .B1(w1[140]), 
        .Y(n21136) );
  AOI22XL U16382 ( .A0(n3028), .A1(w1[20]), .B0(in_valid_w1), .B1(w1[148]), 
        .Y(n21138) );
  AOI222XL U16383 ( .A0(n25567), .A1(w1[33]), .B0(n4576), .B1(w1[1]), .C0(
        w1[129]), .C1(n3216), .Y(n1759) );
  AOI222XL U16384 ( .A0(n25567), .A1(w1[41]), .B0(n4578), .B1(w1[9]), .C0(
        w1[137]), .C1(n3216), .Y(n1791) );
  AOI222XL U16385 ( .A0(n25567), .A1(w1[78]), .B0(n4577), .B1(w1[46]), .C0(
        w1[174]), .C1(n3216), .Y(n1808) );
  AOI222XL U16386 ( .A0(n25567), .A1(w1[108]), .B0(n4577), .B1(w1[76]), .C0(
        w1[204]), .C1(n3216), .Y(n1801) );
  AOI222XL U16387 ( .A0(n25567), .A1(w1[200]), .B0(n3113), .B1(w1[168]), .C0(
        w1[296]), .C1(n3216), .Y(n1912) );
  AOI222XL U16388 ( .A0(n25567), .A1(w1[201]), .B0(n21113), .B1(w1[169]), .C0(
        w1[297]), .C1(n3216), .Y(n1916) );
  AOI222XL U16389 ( .A0(n23088), .A1(w1[202]), .B0(n4577), .B1(w1[170]), .C0(
        w1[298]), .C1(n3216), .Y(n1920) );
  AOI222XL U16390 ( .A0(n25567), .A1(w1[93]), .B0(n3216), .B1(w1[189]), .C0(
        w1[61]), .C1(n25410), .Y(n1868) );
  AOI222XL U16391 ( .A0(n25567), .A1(w1[66]), .B0(n4577), .B1(w1[34]), .C0(
        w1[162]), .C1(n3216), .Y(n1760) );
  AOI222XL U16392 ( .A0(n25567), .A1(w1[67]), .B0(n3113), .B1(w1[35]), .C0(
        w1[163]), .C1(n25541), .Y(n1764) );
  AOI222XL U16393 ( .A0(n25567), .A1(w1[69]), .B0(n4578), .B1(w1[37]), .C0(
        w1[165]), .C1(n25541), .Y(n1772) );
  AOI222XL U16394 ( .A0(n25567), .A1(w1[191]), .B0(n4576), .B1(w1[159]), .C0(
        w1[287]), .C1(n3216), .Y(n2007) );
  AOI222XL U16395 ( .A0(n3061), .A1(w1[106]), .B0(n3051), .B1(w1[74]), .C0(
        w1[202]), .C1(n3216), .Y(n1793) );
  AOI22XL U16396 ( .A0(n3028), .A1(w1[29]), .B0(w1[157]), .B1(in_valid_w1), 
        .Y(n25118) );
  AOI22XL U16397 ( .A0(n3064), .A1(w1[144]), .B0(in_valid_w1), .B1(w1[272]), 
        .Y(n25442) );
  AOI22XL U16398 ( .A0(n3028), .A1(w1[13]), .B0(in_valid_w1), .B1(w1[141]), 
        .Y(n25481) );
  AOI22XL U16399 ( .A0(n3064), .A1(w1[14]), .B0(in_valid_w1), .B1(w1[142]), 
        .Y(n25469) );
  AOI22XL U16400 ( .A0(n3028), .A1(w1[31]), .B0(in_valid_w1), .B1(w1[159]), 
        .Y(n21144) );
  AOI22XL U16401 ( .A0(n3064), .A1(w1[7]), .B0(in_valid_w1), .B1(w1[135]), .Y(
        n21124) );
  AOI22XL U16402 ( .A0(n3028), .A1(w1[9]), .B0(in_valid_w1), .B1(w1[137]), .Y(
        n21128) );
  AOI22XL U16403 ( .A0(n3028), .A1(w1[10]), .B0(in_valid_w1), .B1(w1[138]), 
        .Y(n21150) );
  AOI22XL U16404 ( .A0(n3064), .A1(w1[17]), .B0(in_valid_w1), .B1(w1[145]), 
        .Y(n25432) );
  AOI22XL U16405 ( .A0(n3028), .A1(w1[21]), .B0(in_valid_w1), .B1(w1[149]), 
        .Y(n21140) );
  AOI22XL U16406 ( .A0(n3028), .A1(w1[24]), .B0(w1[152]), .B1(in_valid_w1), 
        .Y(n21142) );
  AOI22XL U16407 ( .A0(n3023), .A1(n26317), .B0(n3061), .B1(n26053), .Y(n25651) );
  AOI22XL U16408 ( .A0(n3023), .A1(n26064), .B0(n25542), .B1(n26360), .Y(
        n25543) );
  AOI22XL U16409 ( .A0(n3023), .A1(n26063), .B0(n25542), .B1(n26359), .Y(
        n25526) );
  AOI22XL U16410 ( .A0(n3023), .A1(n26090), .B0(n3061), .B1(n26392), .Y(n25540) );
  AOI22XL U16411 ( .A0(n3023), .A1(n26089), .B0(n25542), .B1(n26391), .Y(
        n25525) );
  AOI22XL U16412 ( .A0(n3023), .A1(n26057), .B0(n3061), .B1(n26373), .Y(n24372) );
  AOI22XL U16413 ( .A0(n3023), .A1(n26055), .B0(n3061), .B1(n26371), .Y(n24079) );
  AOI22XL U16414 ( .A0(n3023), .A1(n26100), .B0(n3061), .B1(n26355), .Y(n24458) );
  AOI22XL U16415 ( .A0(n3023), .A1(n26079), .B0(n23088), .B1(n26395), .Y(
        n25573) );
  AOI22XL U16416 ( .A0(n3023), .A1(n26069), .B0(n26352), .B1(n3061), .Y(n25087) );
  AOI22XL U16417 ( .A0(n3052), .A1(n26323), .B0(n3061), .B1(n26056), .Y(n25079) );
  AOI22XL U16418 ( .A0(n3052), .A1(n26056), .B0(n3061), .B1(n26374), .Y(n25086) );
  AOI22XL U16419 ( .A0(n3052), .A1(n26101), .B0(n3061), .B1(n26375), .Y(n25114) );
  AOI22XL U16420 ( .A0(n25410), .A1(n26096), .B0(n3061), .B1(n26406), .Y(
        n25574) );
  OAI2BB1XL U16421 ( .A0N(w1[249]), .A1N(n25410), .B0(n24364), .Y(n24365) );
  AOI22XL U16422 ( .A0(n3028), .A1(w1[153]), .B0(w1[281]), .B1(in_valid_w1), 
        .Y(n24364) );
  OAI2BB1XL U16423 ( .A0N(w1[251]), .A1N(n25410), .B0(n25084), .Y(n25085) );
  AOI22XL U16424 ( .A0(n3028), .A1(w1[155]), .B0(w1[283]), .B1(in_valid_w1), 
        .Y(n25084) );
  OAI2BB1XL U16425 ( .A0N(w1[253]), .A1N(n25410), .B0(n25115), .Y(n25116) );
  AOI22XL U16426 ( .A0(n3028), .A1(w1[157]), .B0(w1[285]), .B1(in_valid_w1), 
        .Y(n25115) );
  OAI2BB1XL U16427 ( .A0N(w1[247]), .A1N(n25410), .B0(n24326), .Y(n24327) );
  AOI22XL U16428 ( .A0(n3028), .A1(w1[151]), .B0(w1[279]), .B1(in_valid_w1), 
        .Y(n24326) );
  OAI2BB1XL U16429 ( .A0N(w1[243]), .A1N(n25410), .B0(n25400), .Y(n25401) );
  AOI22XL U16430 ( .A0(n3028), .A1(w1[147]), .B0(in_valid_w1), .B1(w1[275]), 
        .Y(n25400) );
  OAI2BB1XL U16431 ( .A0N(w1[115]), .A1N(n25410), .B0(n25404), .Y(n25405) );
  AOI22XL U16432 ( .A0(n3028), .A1(w1[19]), .B0(in_valid_w1), .B1(w1[147]), 
        .Y(n25404) );
  OAI2BB1XL U16433 ( .A0N(w1[248]), .A1N(n25410), .B0(n21154), .Y(n21155) );
  AOI22XL U16434 ( .A0(n3028), .A1(w1[152]), .B0(w1[280]), .B1(in_valid_w1), 
        .Y(n21154) );
  OAI2BB1XL U16435 ( .A0N(w1[118]), .A1N(n25410), .B0(n21156), .Y(n21157) );
  AOI22XL U16436 ( .A0(n3028), .A1(w1[22]), .B0(in_valid_w1), .B1(w1[150]), 
        .Y(n21156) );
  OAI2BB1XL U16437 ( .A0N(w1[255]), .A1N(n25410), .B0(n21148), .Y(n21149) );
  AOI22XL U16438 ( .A0(n3028), .A1(w1[159]), .B0(in_valid_w1), .B1(w1[287]), 
        .Y(n21148) );
  OAI2BB1XL U16439 ( .A0N(w1[246]), .A1N(n25410), .B0(n21164), .Y(n21165) );
  AOI22XL U16440 ( .A0(n3028), .A1(w1[150]), .B0(in_valid_w1), .B1(w1[278]), 
        .Y(n21164) );
  OAI2BB1XL U16441 ( .A0N(w1[244]), .A1N(n25410), .B0(n21162), .Y(n21163) );
  AOI22XL U16442 ( .A0(n3028), .A1(w1[148]), .B0(in_valid_w1), .B1(w1[276]), 
        .Y(n21162) );
  OAI2BB1XL U16443 ( .A0N(w1[245]), .A1N(n25410), .B0(n21160), .Y(n21161) );
  AOI22XL U16444 ( .A0(n3028), .A1(w1[149]), .B0(in_valid_w1), .B1(w1[277]), 
        .Y(n21160) );
  OAI2BB1XL U16445 ( .A0N(w1[100]), .A1N(n3052), .B0(n25588), .Y(n25589) );
  AOI22XL U16446 ( .A0(n3028), .A1(w1[4]), .B0(in_valid_w1), .B1(w1[132]), .Y(
        n25588) );
  OAI2BB1XL U16447 ( .A0N(w1[227]), .A1N(n3052), .B0(n25603), .Y(n25604) );
  AOI22XL U16448 ( .A0(n3028), .A1(w1[131]), .B0(in_valid_w1), .B1(w1[259]), 
        .Y(n25603) );
  OAI2BB1XL U16449 ( .A0N(w1[102]), .A1N(n3052), .B0(n21146), .Y(n21147) );
  AOI22XL U16450 ( .A0(n3064), .A1(w1[6]), .B0(in_valid_w1), .B1(w1[134]), .Y(
        n21146) );
  OAI2BB1XL U16451 ( .A0N(w1[230]), .A1N(n3052), .B0(n21152), .Y(n21153) );
  AOI22XL U16452 ( .A0(n3064), .A1(w1[134]), .B0(in_valid_w1), .B1(w1[262]), 
        .Y(n21152) );
  OAI2BB1XL U16453 ( .A0N(w1[101]), .A1N(n3052), .B0(n21118), .Y(n21119) );
  AOI22XL U16454 ( .A0(n3064), .A1(w1[5]), .B0(in_valid_w1), .B1(w1[133]), .Y(
        n21118) );
  OAI2BB1XL U16455 ( .A0N(w1[233]), .A1N(n3052), .B0(n21114), .Y(n21115) );
  AOI22XL U16456 ( .A0(n3028), .A1(w1[137]), .B0(in_valid_w1), .B1(w1[265]), 
        .Y(n21114) );
  OAI2BB1XL U16457 ( .A0N(w1[224]), .A1N(n3052), .B0(n25648), .Y(n25649) );
  AOI22XL U16458 ( .A0(n3028), .A1(w1[128]), .B0(in_valid_w1), .B1(w1[256]), 
        .Y(n25648) );
  OAI2BB1XL U16459 ( .A0N(w1[228]), .A1N(n3052), .B0(n25585), .Y(n25586) );
  AOI22XL U16460 ( .A0(n3028), .A1(w1[132]), .B0(in_valid_w1), .B1(w1[260]), 
        .Y(n25585) );
  OAI2BB1XL U16461 ( .A0N(w1[96]), .A1N(n25410), .B0(n25654), .Y(n25655) );
  AOI22XL U16462 ( .A0(n25848), .A1(w1[0]), .B0(in_valid_w1), .B1(w1[128]), 
        .Y(n25654) );
  OAI2BB1XL U16463 ( .A0N(w1[250]), .A1N(n25410), .B0(n24077), .Y(n24078) );
  AOI22XL U16464 ( .A0(n3028), .A1(w1[154]), .B0(w1[282]), .B1(in_valid_w1), 
        .Y(n24077) );
  OAI2BB1XL U16465 ( .A0N(w1[254]), .A1N(n25410), .B0(n25846), .Y(n25847) );
  AOI22XL U16466 ( .A0(n3028), .A1(w1[158]), .B0(w1[286]), .B1(in_valid_w1), 
        .Y(n25846) );
  OAI2BB1XL U16467 ( .A0N(w1[97]), .A1N(n25410), .B0(n25633), .Y(n25634) );
  AOI22XL U16468 ( .A0(n3028), .A1(w1[1]), .B0(in_valid_w1), .B1(w1[129]), .Y(
        n25633) );
  OAI2BB1XL U16469 ( .A0N(w1[225]), .A1N(n25410), .B0(n25630), .Y(n25631) );
  AOI22XL U16470 ( .A0(n3028), .A1(w1[129]), .B0(in_valid_w1), .B1(w1[257]), 
        .Y(n25630) );
  OAI2BB1XL U16471 ( .A0N(w1[226]), .A1N(n25410), .B0(n25617), .Y(n25618) );
  AOI22XL U16472 ( .A0(n3028), .A1(w1[130]), .B0(in_valid_w1), .B1(w1[258]), 
        .Y(n25617) );
  OAI2BB1XL U16473 ( .A0N(w1[114]), .A1N(n25410), .B0(n25418), .Y(n25419) );
  AOI22XL U16474 ( .A0(n3028), .A1(w1[18]), .B0(in_valid_w1), .B1(w1[146]), 
        .Y(n25418) );
  OAI2BB1XL U16475 ( .A0N(w1[237]), .A1N(n25410), .B0(n25479), .Y(n25480) );
  AOI22XL U16476 ( .A0(n3064), .A1(w1[141]), .B0(in_valid_w1), .B1(w1[269]), 
        .Y(n25479) );
  OAI2BB1XL U16477 ( .A0N(w1[238]), .A1N(n25410), .B0(n25466), .Y(n25467) );
  AOI22XL U16478 ( .A0(n3064), .A1(w1[142]), .B0(in_valid_w1), .B1(w1[270]), 
        .Y(n25466) );
  OAI2BB1XL U16479 ( .A0N(w1[239]), .A1N(n25410), .B0(n25454), .Y(n25455) );
  AOI22XL U16480 ( .A0(n3064), .A1(w1[143]), .B0(in_valid_w1), .B1(w1[271]), 
        .Y(n25454) );
  OAI2BB1XL U16481 ( .A0N(w1[241]), .A1N(n25410), .B0(n25429), .Y(n25430) );
  AOI22XL U16482 ( .A0(n3064), .A1(w1[145]), .B0(in_valid_w1), .B1(w1[273]), 
        .Y(n25429) );
  OAI2BB1XL U16483 ( .A0N(w1[242]), .A1N(n25410), .B0(n25415), .Y(n25416) );
  AOI22XL U16484 ( .A0(n3028), .A1(w1[146]), .B0(in_valid_w1), .B1(w1[274]), 
        .Y(n25415) );
  OAI2BB1XL U16485 ( .A0N(w1[229]), .A1N(n25410), .B0(n21130), .Y(n21131) );
  AOI22XL U16486 ( .A0(n3064), .A1(w1[133]), .B0(in_valid_w1), .B1(w1[261]), 
        .Y(n21130) );
  OAI2BB1XL U16487 ( .A0N(w1[231]), .A1N(n25410), .B0(n21120), .Y(n21121) );
  AOI22XL U16488 ( .A0(n3064), .A1(w1[135]), .B0(in_valid_w1), .B1(w1[263]), 
        .Y(n21120) );
  OAI2BB1XL U16489 ( .A0N(w1[235]), .A1N(n25410), .B0(n21158), .Y(n21159) );
  AOI22XL U16490 ( .A0(n3064), .A1(w1[139]), .B0(in_valid_w1), .B1(w1[267]), 
        .Y(n21158) );
  OAI2BB1XL U16491 ( .A0N(w1[236]), .A1N(n25410), .B0(n21134), .Y(n21135) );
  AOI22XL U16492 ( .A0(n3028), .A1(w1[140]), .B0(in_valid_w1), .B1(w1[268]), 
        .Y(n21134) );
  OAI2BB1XL U16493 ( .A0N(w1[232]), .A1N(n25410), .B0(n21122), .Y(n21123) );
  AOI22XL U16494 ( .A0(n3064), .A1(w1[136]), .B0(in_valid_w1), .B1(w1[264]), 
        .Y(n21122) );
  OAI2BB1XL U16495 ( .A0N(w1[234]), .A1N(n25410), .B0(n21116), .Y(n21117) );
  AOI22XL U16496 ( .A0(n3028), .A1(w1[138]), .B0(in_valid_w1), .B1(w1[266]), 
        .Y(n21116) );
  AOI22XL U16497 ( .A0(n3052), .A1(n26071), .B0(n25542), .B1(n26364), .Y(
        n25431) );
  AOI22XL U16498 ( .A0(n3052), .A1(n26325), .B0(n3061), .B1(n26059), .Y(n25802) );
  AOI22XL U16499 ( .A0(n3052), .A1(n26094), .B0(n3061), .B1(n26404), .Y(n25417) );
  AOI22XL U16500 ( .A0(n3052), .A1(n26084), .B0(n3061), .B1(n26384), .Y(n25427) );
  AOI22XL U16501 ( .A0(n3052), .A1(n26050), .B0(n23088), .B1(n26383), .Y(
        n25413) );
  AOI22XL U16502 ( .A0(n3052), .A1(n26104), .B0(n3061), .B1(n26361), .Y(n25444) );
  AOI22XL U16503 ( .A0(n3052), .A1(n26054), .B0(n3061), .B1(n26403), .Y(n25402) );
  AOI22XL U16504 ( .A0(n3052), .A1(n26077), .B0(n3061), .B1(n26382), .Y(n25398) );
  AOI22XL U16505 ( .A0(n3052), .A1(n26083), .B0(n3061), .B1(n26381), .Y(n25390) );
  AOI22XL U16506 ( .A0(n3052), .A1(n26065), .B0(n3061), .B1(n26356), .Y(n25399) );
  AOI22XL U16507 ( .A0(n3052), .A1(n26326), .B0(n3061), .B1(n26054), .Y(n25403) );
  AOI222XL U16508 ( .A0(n25567), .A1(w1[91]), .B0(n3216), .B1(w1[187]), .C0(
        w1[59]), .C1(n25410), .Y(n1860) );
  AOI22XL U16509 ( .A0(n3052), .A1(n26322), .B0(n3061), .B1(n26055), .Y(n24080) );
  AOI22XL U16510 ( .A0(n3052), .A1(n26099), .B0(n3061), .B1(n26372), .Y(n24322) );
  AOI22XL U16511 ( .A0(n3052), .A1(n26319), .B0(n3061), .B1(n26050), .Y(n25414) );
  AOI22XL U16512 ( .A0(n3052), .A1(n26066), .B0(n3061), .B1(n26357), .Y(n25441) );
  AOI22XL U16513 ( .A0(n3052), .A1(n26074), .B0(n25542), .B1(n26388), .Y(
        n25491) );
  AOI22XL U16514 ( .A0(n3052), .A1(n26098), .B0(n25542), .B1(n26408), .Y(
        n25632) );
  AOI22XL U16515 ( .A0(n3064), .A1(w1[15]), .B0(in_valid_w1), .B1(w1[143]), 
        .Y(n25456) );
  AOI22XL U16516 ( .A0(n3064), .A1(w1[16]), .B0(in_valid_w1), .B1(w1[144]), 
        .Y(n25445) );
  AOI22XL U16517 ( .A0(n25410), .A1(n26062), .B0(n3061), .B1(n26358), .Y(
        n25515) );
  AOI22XL U16518 ( .A0(n25410), .A1(n26082), .B0(n3061), .B1(n26380), .Y(
        n25377) );
  AOI22XL U16519 ( .A0(n3023), .A1(n26076), .B0(n3061), .B1(n26379), .Y(n25368) );
  AOI22XL U16520 ( .A0(n25410), .A1(n26093), .B0(n3061), .B1(n26402), .Y(
        n25369) );
  AOI22XL U16521 ( .A0(n3028), .A1(w1[25]), .B0(w1[153]), .B1(in_valid_w1), 
        .Y(n24366) );
  AOI22XL U16522 ( .A0(n3028), .A1(w1[28]), .B0(w1[156]), .B1(in_valid_w1), 
        .Y(n24452) );
  AOI22XL U16523 ( .A0(n25848), .A1(w1[30]), .B0(w1[158]), .B1(in_valid_w1), 
        .Y(n25849) );
  AOI22XL U16524 ( .A0(n3028), .A1(w1[23]), .B0(w1[151]), .B1(in_valid_w1), 
        .Y(n24328) );
  AOI22XL U16525 ( .A0(n3028), .A1(w1[26]), .B0(w1[154]), .B1(in_valid_w1), 
        .Y(n24081) );
  MXI2X1 U16526 ( .A(data[46]), .B(data[78]), .S0(n3229), .Y(n1660) );
  MXI2XL U16527 ( .A(data[47]), .B(data[79]), .S0(n3229), .Y(n1661) );
  MXI2XL U16528 ( .A(data[48]), .B(data[80]), .S0(n3123), .Y(n1662) );
  MXI2XL U16529 ( .A(data[50]), .B(data[82]), .S0(n3229), .Y(n1664) );
  MXI2XL U16530 ( .A(data[76]), .B(data[108]), .S0(n3123), .Y(n1690) );
  MXI2XL U16531 ( .A(data[83]), .B(data[115]), .S0(n3229), .Y(n1697) );
  MXI2XL U16532 ( .A(data[35]), .B(data[67]), .S0(n3229), .Y(n1649) );
  MXI2XL U16533 ( .A(data[37]), .B(data[69]), .S0(n3229), .Y(n1651) );
  MXI2XL U16534 ( .A(data[38]), .B(data[70]), .S0(n3123), .Y(n1652) );
  MXI2XL U16535 ( .A(data[39]), .B(data[71]), .S0(n3229), .Y(n1653) );
  MXI2XL U16536 ( .A(data[40]), .B(data[72]), .S0(n3229), .Y(n1654) );
  MXI2XL U16537 ( .A(data[41]), .B(data[73]), .S0(n3229), .Y(n1655) );
  MXI2XL U16538 ( .A(data[42]), .B(data[74]), .S0(n3229), .Y(n1656) );
  MXI2XL U16539 ( .A(data[43]), .B(data[75]), .S0(n3123), .Y(n1657) );
  MXI2XL U16540 ( .A(data[44]), .B(data[76]), .S0(n3229), .Y(n1658) );
  MXI2XL U16541 ( .A(data[49]), .B(data[81]), .S0(n3123), .Y(n1663) );
  MXI2XL U16542 ( .A(data[52]), .B(data[84]), .S0(n3123), .Y(n1666) );
  MXI2XL U16543 ( .A(data[53]), .B(data[85]), .S0(n3229), .Y(n1667) );
  MXI2XL U16544 ( .A(data[54]), .B(data[86]), .S0(n3123), .Y(n1668) );
  MXI2XL U16545 ( .A(data[70]), .B(data[102]), .S0(n3123), .Y(n1684) );
  MXI2XL U16546 ( .A(data[71]), .B(data[103]), .S0(n4579), .Y(n1685) );
  MXI2XL U16547 ( .A(data[72]), .B(data[104]), .S0(n4579), .Y(n1686) );
  MXI2XL U16548 ( .A(data[73]), .B(data[105]), .S0(n3229), .Y(n1687) );
  MXI2XL U16549 ( .A(data[74]), .B(data[106]), .S0(n4579), .Y(n1688) );
  MXI2XL U16550 ( .A(data[75]), .B(data[107]), .S0(n4579), .Y(n1689) );
  MXI2XL U16551 ( .A(data[78]), .B(data[110]), .S0(n4579), .Y(n1692) );
  MXI2XL U16552 ( .A(data[79]), .B(data[111]), .S0(n4579), .Y(n1693) );
  MXI2XL U16553 ( .A(data[80]), .B(data[112]), .S0(n4579), .Y(n1694) );
  MXI2XL U16554 ( .A(data[81]), .B(data[113]), .S0(n4579), .Y(n1695) );
  MXI2XL U16555 ( .A(data[82]), .B(data[114]), .S0(n4579), .Y(n1696) );
  MXI2XL U16556 ( .A(data[84]), .B(data[116]), .S0(n4579), .Y(n1698) );
  MXI2XL U16557 ( .A(data[85]), .B(data[117]), .S0(n4579), .Y(n1699) );
  MXI2XL U16558 ( .A(data[32]), .B(data[64]), .S0(n3123), .Y(n1646) );
  MXI2XL U16559 ( .A(data[33]), .B(data[65]), .S0(n3123), .Y(n1647) );
  MXI2XL U16560 ( .A(data[34]), .B(data[66]), .S0(n3123), .Y(n1648) );
  MXI2XL U16561 ( .A(data[36]), .B(data[68]), .S0(n3123), .Y(n1650) );
  MXI2XL U16562 ( .A(data[45]), .B(data[77]), .S0(n3123), .Y(n1659) );
  MXI2XL U16563 ( .A(data[51]), .B(data[83]), .S0(n3123), .Y(n1665) );
  MXI2XL U16564 ( .A(data[64]), .B(data[96]), .S0(n3123), .Y(n1678) );
  MXI2XL U16565 ( .A(data[65]), .B(data[97]), .S0(n3229), .Y(n1679) );
  MXI2XL U16566 ( .A(data[66]), .B(data[98]), .S0(n3229), .Y(n1680) );
  MXI2XL U16567 ( .A(data[67]), .B(data[99]), .S0(n3229), .Y(n1681) );
  MXI2XL U16568 ( .A(data[68]), .B(data[100]), .S0(n3229), .Y(n1682) );
  MXI2XL U16569 ( .A(data[69]), .B(data[101]), .S0(n3229), .Y(n1683) );
  MXI2XL U16570 ( .A(data[77]), .B(data[109]), .S0(n3229), .Y(n1691) );
  MXI2XL U16571 ( .A(data[86]), .B(data[118]), .S0(n3229), .Y(n1700) );
  AOI22XL U16572 ( .A0(n24739), .A1(y10[26]), .B0(n3050), .B1(y12[26]), .Y(
        n24418) );
  AOI22XL U16573 ( .A0(n24739), .A1(y10[30]), .B0(n3050), .B1(y12[30]), .Y(
        n23694) );
  AOI22XL U16574 ( .A0(n24739), .A1(y10[11]), .B0(n25656), .B1(y12[11]), .Y(
        n23655) );
  AOI22XL U16575 ( .A0(n24739), .A1(y10[10]), .B0(n8104), .B1(y12[10]), .Y(
        n24641) );
  AOI22XL U16576 ( .A0(n24739), .A1(y10[9]), .B0(n25656), .B1(y12[9]), .Y(
        n23576) );
  AOI22XL U16577 ( .A0(n24739), .A1(y10[4]), .B0(n25656), .B1(y12[4]), .Y(
        n24522) );
  AOI22XL U16578 ( .A0(n25025), .A1(y10[16]), .B0(n25656), .B1(y12[16]), .Y(
        n23755) );
  AOI22XL U16579 ( .A0(n24739), .A1(y10[13]), .B0(n25656), .B1(y12[13]), .Y(
        n24713) );
  NAND2XL U16580 ( .A(in_valid_w2), .B(weight2[1]), .Y(n25032) );
  AOI2BB1XL U16581 ( .A0N(n25611), .A1N(n3118), .B0(n25068), .Y(n2202) );
  NAND2XL U16582 ( .A(in_valid_w2), .B(weight2[2]), .Y(n25067) );
  NAND2XL U16583 ( .A(in_valid_w2), .B(weight2[3]), .Y(n25034) );
  AOI2BB1XL U16584 ( .A0N(n25579), .A1N(n3118), .B0(n25066), .Y(n2204) );
  NAND2XL U16585 ( .A(in_valid_w2), .B(weight2[4]), .Y(n25065) );
  NAND2XL U16586 ( .A(in_valid_w2), .B(weight2[5]), .Y(n25036) );
  AOI2BB1XL U16587 ( .A0N(n25559), .A1N(n3118), .B0(n25064), .Y(n2206) );
  NAND2XL U16588 ( .A(in_valid_w2), .B(weight2[6]), .Y(n25063) );
  NAND2XL U16589 ( .A(in_valid_w2), .B(weight2[7]), .Y(n25038) );
  AOI2BB1XL U16590 ( .A0N(n25536), .A1N(n3118), .B0(n25062), .Y(n2208) );
  NAND2XL U16591 ( .A(in_valid_w2), .B(weight2[8]), .Y(n25061) );
  NAND2XL U16592 ( .A(in_valid_w2), .B(weight2[9]), .Y(n25040) );
  AOI2BB1XL U16593 ( .A0N(n25510), .A1N(n3118), .B0(n25060), .Y(n2210) );
  NAND2XL U16594 ( .A(in_valid_w2), .B(weight2[10]), .Y(n25058) );
  NAND2XL U16595 ( .A(in_valid_w2), .B(weight2[11]), .Y(n25042) );
  AOI2BB1XL U16596 ( .A0N(n25487), .A1N(n3118), .B0(n25057), .Y(n2212) );
  NAND2XL U16597 ( .A(in_valid_w2), .B(weight2[12]), .Y(n25056) );
  NAND2XL U16598 ( .A(in_valid_w2), .B(weight2[13]), .Y(n25044) );
  NAND2XL U16599 ( .A(in_valid_w2), .B(weight2[14]), .Y(n15907) );
  AOI2BB1XL U16600 ( .A0N(n25449), .A1N(n3118), .B0(n25047), .Y(n2215) );
  NAND2XL U16601 ( .A(in_valid_w2), .B(weight2[15]), .Y(n25046) );
  NAND2XL U16602 ( .A(in_valid_w2), .B(weight2[16]), .Y(n15938) );
  NAND2XL U16603 ( .A(in_valid_w2), .B(weight2[17]), .Y(n21015) );
  AOI2BB1XL U16604 ( .A0N(n25408), .A1N(n3118), .B0(n25055), .Y(n2218) );
  NAND2XL U16605 ( .A(in_valid_w2), .B(weight2[18]), .Y(n25054) );
  AOI2BB1XL U16606 ( .A0N(n25394), .A1N(n3118), .B0(n25049), .Y(n2219) );
  NAND2XL U16607 ( .A(in_valid_w2), .B(weight2[19]), .Y(n25048) );
  AOI2BB1XL U16608 ( .A0N(n25386), .A1N(n3118), .B0(n25053), .Y(n2220) );
  NAND2XL U16609 ( .A(in_valid_w2), .B(weight2[20]), .Y(n25052) );
  AOI2BB1XL U16610 ( .A0N(n25373), .A1N(n3118), .B0(n25051), .Y(n2221) );
  NAND2XL U16611 ( .A(in_valid_w2), .B(weight2[21]), .Y(n25050) );
  OAI21XL U16612 ( .A0(n24421), .A1(n25711), .B0(n23814), .Y(n2161) );
  AOI22XL U16613 ( .A0(n25820), .A1(n26042), .B0(in_valid_w2), .B1(n26423), 
        .Y(n23814) );
  OAI21XL U16614 ( .A0(n24417), .A1(n25711), .B0(n23820), .Y(n2162) );
  AOI22XL U16615 ( .A0(n25822), .A1(n26043), .B0(in_valid_w2), .B1(n26298), 
        .Y(n23820) );
  OAI21XL U16616 ( .A0(n25080), .A1(n25711), .B0(n25078), .Y(n2163) );
  AOI22XL U16617 ( .A0(n25822), .A1(n26045), .B0(in_valid_w2), .B1(n26421), 
        .Y(n25078) );
  OAI21XL U16618 ( .A0(n24451), .A1(n25711), .B0(n24450), .Y(n2164) );
  AOI22XL U16619 ( .A0(n25822), .A1(n26301), .B0(in_valid_w2), .B1(n26044), 
        .Y(n24450) );
  OAI21XL U16620 ( .A0(n25683), .A1(n25711), .B0(n23848), .Y(n2165) );
  AOI22XL U16621 ( .A0(n25822), .A1(n26047), .B0(in_valid_w2), .B1(n26422), 
        .Y(n23848) );
  OAI21XL U16622 ( .A0(n25801), .A1(n25711), .B0(n23838), .Y(n2166) );
  AOI22XL U16623 ( .A0(n25822), .A1(n26046), .B0(in_valid_w2), .B1(n26304), 
        .Y(n23838) );
  OAI21XL U16624 ( .A0(n24769), .A1(n3059), .B0(n24766), .Y(n24767) );
  OAI21XL U16625 ( .A0(n24821), .A1(n3059), .B0(n24818), .Y(n24819) );
  OAI21XL U16626 ( .A0(n24321), .A1(n25711), .B0(n23971), .Y(n2159) );
  AOI22XL U16627 ( .A0(n25820), .A1(n26037), .B0(in_valid_w2), .B1(n26285), 
        .Y(n23971) );
  AOI22XL U16628 ( .A0(n25820), .A1(n26036), .B0(in_valid_w2), .B1(n26284), 
        .Y(n25710) );
  AOI21XL U16629 ( .A0(n24510), .A1(n24525), .B0(n24509), .Y(n2399) );
  AOI22XL U16630 ( .A0(n24958), .A1(y12[3]), .B0(n3050), .B1(y11[3]), .Y(
        n24508) );
  AOI22XL U16631 ( .A0(n25815), .A1(y12[7]), .B0(n25656), .B1(y11[7]), .Y(
        n24592) );
  AOI22XL U16632 ( .A0(n25815), .A1(y12[8]), .B0(n25656), .B1(y11[8]), .Y(
        n24604) );
  AOI21XL U16633 ( .A0(n24738), .A1(n3060), .B0(n24737), .Y(n2421) );
  INVXL U16634 ( .A(n24735), .Y(n24738) );
  AOI22XL U16635 ( .A0(n24739), .A1(y12[14]), .B0(n8104), .B1(y11[14]), .Y(
        n24736) );
  AOI21XL U16636 ( .A0(n24887), .A1(n6161), .B0(n24886), .Y(n2429) );
  AOI22XL U16637 ( .A0(n25025), .A1(y12[18]), .B0(n3050), .B1(y11[18]), .Y(
        n24885) );
  AOI21XL U16638 ( .A0(n24983), .A1(n3060), .B0(n24982), .Y(n2433) );
  AOI22XL U16639 ( .A0(n25025), .A1(y12[20]), .B0(n3050), .B1(y11[20]), .Y(
        n24981) );
  AOI22XL U16640 ( .A0(n25025), .A1(y12[21]), .B0(n3050), .B1(y11[21]), .Y(
        n25026) );
  AOI21XL U16641 ( .A0(n25339), .A1(n6161), .B0(n25338), .Y(n2437) );
  AOI22XL U16642 ( .A0(n24958), .A1(y12[23]), .B0(n3050), .B1(y11[23]), .Y(
        n24316) );
  NOR2X1 U16643 ( .A(n5085), .B(n25693), .Y(n5084) );
  NAND2X1 U16644 ( .A(n19089), .B(n3120), .Y(n4936) );
  OAI21XL U16645 ( .A0(n24149), .A1(n25328), .B0(n5311), .Y(n5310) );
  AOI22XL U16646 ( .A0(n22486), .A1(sigma11[0]), .B0(n25754), .B1(sigma12[0]), 
        .Y(n25332) );
  NOR2X1 U16647 ( .A(n5085), .B(n25255), .Y(n24056) );
  AOI22XL U16648 ( .A0(n22486), .A1(sigma12[1]), .B0(n25750), .B1(sigma11[1]), 
        .Y(n24054) );
  AOI22XL U16649 ( .A0(n22486), .A1(sigma12[6]), .B0(n25750), .B1(sigma11[6]), 
        .Y(n24141) );
  NAND2X1 U16650 ( .A(n5879), .B(n24196), .Y(n24197) );
  AOI22XL U16651 ( .A0(n22486), .A1(sigma12[14]), .B0(n25750), .B1(sigma11[14]), .Y(n24196) );
  AOI22XL U16652 ( .A0(n22486), .A1(sigma12[18]), .B0(n25750), .B1(sigma11[18]), .Y(n24232) );
  AOI22XL U16653 ( .A0(n22486), .A1(sigma11[13]), .B0(n25754), .B1(sigma12[13]), .Y(n24193) );
  AOI22XL U16654 ( .A0(n22486), .A1(sigma12[5]), .B0(n25750), .B1(sigma11[5]), 
        .Y(n24131) );
  AOI22XL U16655 ( .A0(n22486), .A1(sigma12[8]), .B0(n25750), .B1(sigma11[8]), 
        .Y(n24152) );
  AOI22XL U16656 ( .A0(n22486), .A1(sigma12[10]), .B0(n25750), .B1(sigma11[10]), .Y(n24164) );
  AOI22XL U16657 ( .A0(n22486), .A1(sigma12[11]), .B0(n25750), .B1(sigma11[11]), .Y(n24175) );
  AOI22XL U16658 ( .A0(n22486), .A1(sigma12[12]), .B0(n25750), .B1(sigma11[12]), .Y(n24180) );
  AOI211XL U16659 ( .A0(n25761), .A1(n24218), .B0(n24217), .C0(n24216), .Y(
        n2329) );
  OAI21XL U16660 ( .A0(mul5_out[11]), .A1(n4875), .B0(n24176), .Y(n2318) );
  AOI22XL U16661 ( .A0(n25763), .A1(n26517), .B0(n25754), .B1(n26447), .Y(
        n24176) );
  AOI22XL U16662 ( .A0(n25754), .A1(sigma11[7]), .B0(sigma12[7]), .B1(n20748), 
        .Y(n20743) );
  INVXL U16663 ( .A(n20362), .Y(n5948) );
  AOI22XL U16664 ( .A0(n25255), .A1(sigma12[15]), .B0(n3050), .B1(sigma11[15]), 
        .Y(n20362) );
  INVXL U16665 ( .A(n20354), .Y(n5849) );
  AOI22XL U16666 ( .A0(n25754), .A1(sigma11[17]), .B0(sigma12[17]), .B1(n3059), 
        .Y(n20354) );
  AOI22XL U16667 ( .A0(n25255), .A1(sigma12[18]), .B0(n3050), .B1(sigma11[18]), 
        .Y(n21050) );
  AOI22XL U16668 ( .A0(n25255), .A1(sigma12[20]), .B0(n3050), .B1(sigma11[20]), 
        .Y(n20925) );
  AOI22XL U16669 ( .A0(n22486), .A1(sigma11[9]), .B0(n25754), .B1(sigma12[9]), 
        .Y(n24161) );
  AOI22XL U16670 ( .A0(n25754), .A1(sigma11[1]), .B0(sigma12[1]), .B1(n3024), 
        .Y(n20696) );
  NAND2X1 U16671 ( .A(n23697), .B(n25767), .Y(n4852) );
  AOI22XL U16672 ( .A0(n25754), .A1(sigma11[6]), .B0(sigma12[6]), .B1(n3024), 
        .Y(n20937) );
  AOI22XL U16673 ( .A0(n22486), .A1(sigma12[3]), .B0(n25750), .B1(sigma11[3]), 
        .Y(n24118) );
  NOR2X1 U16674 ( .A(n24888), .B(n25255), .Y(n24243) );
  NAND2X1 U16675 ( .A(n5427), .B(n24241), .Y(n24242) );
  AOI22XL U16676 ( .A0(n22486), .A1(sigma12[2]), .B0(n25750), .B1(sigma11[2]), 
        .Y(n24114) );
  OAI21XL U16677 ( .A0(mul5_out[13]), .A1(n5032), .B0(n24191), .Y(n2322) );
  AOI22XL U16678 ( .A0(n25763), .A1(n26032), .B0(n25754), .B1(n26443), .Y(
        n24191) );
  OAI21XL U16679 ( .A0(n24129), .A1(n5032), .B0(n24128), .Y(n24130) );
  AOI22XL U16680 ( .A0(n22486), .A1(sigma12[4]), .B0(n25750), .B1(sigma11[4]), 
        .Y(n24128) );
  AOI22XL U16681 ( .A0(n22486), .A1(sigma12[22]), .B0(n25750), .B1(sigma11[22]), .Y(n25756) );
  AOI22XL U16682 ( .A0(n22486), .A1(sigma12[23]), .B0(n25750), .B1(sigma11[23]), .Y(n25771) );
  AOI22XL U16683 ( .A0(n22486), .A1(sigma12[24]), .B0(n25750), .B1(sigma11[24]), .Y(n25196) );
  OAI21XL U16684 ( .A0(mul5_out[10]), .A1(n4875), .B0(n24168), .Y(n2316) );
  AOI22XL U16685 ( .A0(n25763), .A1(n26516), .B0(n25754), .B1(n26446), .Y(
        n24168) );
  OAI21XL U16686 ( .A0(mul5_out[4]), .A1(n5032), .B0(n20345), .Y(n2304) );
  AOI22XL U16687 ( .A0(n25786), .A1(n26370), .B0(n25785), .B1(n26041), .Y(
        n20345) );
  OAI21XL U16688 ( .A0(n25189), .A1(n5015), .B0(n25188), .Y(n25190) );
  AOI22XL U16689 ( .A0(n22486), .A1(sigma12[25]), .B0(n25750), .B1(sigma11[25]), .Y(n25188) );
  AOI22XL U16690 ( .A0(n25201), .A1(sigma12[26]), .B0(n25750), .B1(sigma11[26]), .Y(n25175) );
  NAND2X1 U16691 ( .A(n6021), .B(n24112), .Y(n24113) );
  AOI21XL U16692 ( .A0(n25754), .A1(n25674), .B0(n25208), .Y(n2355) );
  AOI22XL U16693 ( .A0(n22486), .A1(sigma12[29]), .B0(n17459), .B1(sigma11[29]), .Y(n25205) );
  OAI21XL U16694 ( .A0(n25783), .A1(n5032), .B0(n25782), .Y(n25784) );
  AOI22XL U16695 ( .A0(n22486), .A1(sigma12[30]), .B0(n25750), .B1(sigma11[30]), .Y(n25782) );
  AOI22XL U16696 ( .A0(n3028), .A1(w1[283]), .B0(in_valid_w1), .B1(weight1[27]), .Y(n25081) );
  OAI2BB1XL U16697 ( .A0N(w1[380]), .A1N(n25410), .B0(n24454), .Y(n24455) );
  AOI22XL U16698 ( .A0(n3028), .A1(w1[284]), .B0(in_valid_w1), .B1(weight1[28]), .Y(n24454) );
  OAI21XL U16699 ( .A0(n25533), .A1(n3226), .B0(n25532), .Y(n2041) );
  AOI22XL U16700 ( .A0(n3052), .A1(n26061), .B0(n3061), .B1(n26476), .Y(n25532) );
  OAI21XL U16701 ( .A0(n25518), .A1(n3226), .B0(n25517), .Y(n2045) );
  AOI22XL U16702 ( .A0(n3052), .A1(n26060), .B0(n3061), .B1(n26475), .Y(n25517) );
  OAI21XL U16703 ( .A0(n25677), .A1(n4572), .B0(n25676), .Y(n2009) );
  AOI22XL U16704 ( .A0(n3052), .A1(n26133), .B0(n3061), .B1(n26484), .Y(n25676) );
  OAI21XL U16705 ( .A0(n25623), .A1(n4573), .B0(n25622), .Y(n2013) );
  AOI22XL U16706 ( .A0(n25410), .A1(n26132), .B0(n3061), .B1(n26483), .Y(
        n25622) );
  OAI21XL U16707 ( .A0(n25609), .A1(n3226), .B0(n25608), .Y(n2017) );
  AOI22XL U16708 ( .A0(n3052), .A1(n26131), .B0(n23088), .B1(n26482), .Y(
        n25608) );
  OAI21XL U16709 ( .A0(n25596), .A1(n3226), .B0(n25595), .Y(n2021) );
  AOI22XL U16710 ( .A0(n25410), .A1(n26130), .B0(n3061), .B1(n26481), .Y(
        n25595) );
  OAI21XL U16711 ( .A0(n25495), .A1(n4573), .B0(n25494), .Y(n2053) );
  AOI22XL U16712 ( .A0(n3052), .A1(n26124), .B0(n3061), .B1(n26473), .Y(n25494) );
  OAI21XL U16713 ( .A0(n25472), .A1(n4574), .B0(n25471), .Y(n2061) );
  AOI22XL U16714 ( .A0(n3052), .A1(n26123), .B0(n3061), .B1(n26471), .Y(n25471) );
  OAI21XL U16715 ( .A0(n25448), .A1(n4572), .B0(n25447), .Y(n2069) );
  AOI22XL U16716 ( .A0(n3052), .A1(n26121), .B0(n3061), .B1(n26469), .Y(n25447) );
  OAI21XL U16717 ( .A0(n25421), .A1(n4571), .B0(n25420), .Y(n2077) );
  AOI22XL U16718 ( .A0(n25410), .A1(n26120), .B0(n3061), .B1(n26467), .Y(
        n25420) );
  OAI21XL U16719 ( .A0(n25407), .A1(n4571), .B0(n25406), .Y(n2081) );
  AOI22XL U16720 ( .A0(n3052), .A1(n26119), .B0(n3061), .B1(n26466), .Y(n25406) );
  OAI21XL U16721 ( .A0(n25392), .A1(n25584), .B0(n25391), .Y(n2085) );
  AOI22XL U16722 ( .A0(n3052), .A1(n26118), .B0(n3061), .B1(n26465), .Y(n25391) );
  OAI21XL U16723 ( .A0(n25384), .A1(n25584), .B0(n25383), .Y(n2089) );
  AOI22XL U16724 ( .A0(n3052), .A1(n26117), .B0(n3061), .B1(n26464), .Y(n25383) );
  OAI21XL U16725 ( .A0(n25821), .A1(n25584), .B0(n25364), .Y(n2097) );
  AOI22XL U16726 ( .A0(n3052), .A1(n26115), .B0(n3061), .B1(n26462), .Y(n25364) );
  OAI2BB1XL U16727 ( .A0N(w1[353]), .A1N(n25410), .B0(n25626), .Y(n25627) );
  AOI22XL U16728 ( .A0(n3028), .A1(w1[257]), .B0(in_valid_w1), .B1(weight1[1]), 
        .Y(n25626) );
  OAI2BB1XL U16729 ( .A0N(w1[354]), .A1N(n25410), .B0(n25612), .Y(n25613) );
  AOI22XL U16730 ( .A0(n3028), .A1(w1[258]), .B0(in_valid_w1), .B1(weight1[2]), 
        .Y(n25612) );
  OAI2BB1XL U16731 ( .A0N(w1[355]), .A1N(n3052), .B0(n25599), .Y(n25600) );
  AOI22XL U16732 ( .A0(n3028), .A1(w1[259]), .B0(in_valid_w1), .B1(weight1[3]), 
        .Y(n25599) );
  OAI2BB1XL U16733 ( .A0N(w1[357]), .A1N(n3052), .B0(n25570), .Y(n25571) );
  AOI22XL U16734 ( .A0(n3064), .A1(w1[261]), .B0(in_valid_w1), .B1(weight1[5]), 
        .Y(n25570) );
  OAI2BB1XL U16735 ( .A0N(w1[358]), .A1N(n25410), .B0(n25560), .Y(n25561) );
  AOI22XL U16736 ( .A0(n3064), .A1(w1[262]), .B0(in_valid_w1), .B1(weight1[6]), 
        .Y(n25560) );
  OAI2BB1XL U16737 ( .A0N(w1[359]), .A1N(n3052), .B0(n25548), .Y(n25549) );
  AOI22XL U16738 ( .A0(n3064), .A1(w1[263]), .B0(in_valid_w1), .B1(weight1[7]), 
        .Y(n25548) );
  OAI2BB1XL U16739 ( .A0N(w1[360]), .A1N(n3052), .B0(n25537), .Y(n25538) );
  AOI22XL U16740 ( .A0(n3064), .A1(w1[264]), .B0(in_valid_w1), .B1(weight1[8]), 
        .Y(n25537) );
  OAI2BB1XL U16741 ( .A0N(w1[361]), .A1N(n3052), .B0(n25522), .Y(n25523) );
  AOI22XL U16742 ( .A0(n3064), .A1(w1[265]), .B0(in_valid_w1), .B1(weight1[9]), 
        .Y(n25522) );
  OAI2BB1XL U16743 ( .A0N(w1[362]), .A1N(n25410), .B0(n25511), .Y(n25512) );
  AOI22XL U16744 ( .A0(n3028), .A1(w1[266]), .B0(in_valid_w1), .B1(weight1[10]), .Y(n25511) );
  OAI2BB1XL U16745 ( .A0N(w1[363]), .A1N(n25410), .B0(n25498), .Y(n25499) );
  AOI22XL U16746 ( .A0(n3028), .A1(w1[267]), .B0(in_valid_w1), .B1(weight1[11]), .Y(n25498) );
  OAI2BB1XL U16747 ( .A0N(w1[364]), .A1N(n25410), .B0(n25488), .Y(n25489) );
  AOI22XL U16748 ( .A0(n3064), .A1(w1[268]), .B0(in_valid_w1), .B1(weight1[12]), .Y(n25488) );
  OAI2BB1XL U16749 ( .A0N(w1[365]), .A1N(n3052), .B0(n25474), .Y(n25475) );
  AOI22XL U16750 ( .A0(n3064), .A1(w1[269]), .B0(in_valid_w1), .B1(weight1[13]), .Y(n25474) );
  OAI2BB1XL U16751 ( .A0N(w1[366]), .A1N(n25410), .B0(n25462), .Y(n25463) );
  AOI22XL U16752 ( .A0(n3064), .A1(w1[270]), .B0(in_valid_w1), .B1(weight1[14]), .Y(n25462) );
  OAI2BB1XL U16753 ( .A0N(w1[367]), .A1N(n25410), .B0(n25450), .Y(n25451) );
  AOI22XL U16754 ( .A0(n3064), .A1(w1[271]), .B0(in_valid_w1), .B1(weight1[15]), .Y(n25450) );
  OAI2BB1XL U16755 ( .A0N(w1[368]), .A1N(n3052), .B0(n25438), .Y(n25439) );
  AOI22XL U16756 ( .A0(n3064), .A1(w1[272]), .B0(in_valid_w1), .B1(weight1[16]), .Y(n25438) );
  OAI2BB1XL U16757 ( .A0N(w1[369]), .A1N(n3052), .B0(n25424), .Y(n25425) );
  AOI22XL U16758 ( .A0(n3028), .A1(w1[273]), .B0(in_valid_w1), .B1(weight1[17]), .Y(n25424) );
  OAI2BB1XL U16759 ( .A0N(w1[370]), .A1N(n25410), .B0(n25409), .Y(n25411) );
  AOI22XL U16760 ( .A0(n3028), .A1(w1[274]), .B0(in_valid_w1), .B1(weight1[18]), .Y(n25409) );
  OAI2BB1XL U16761 ( .A0N(w1[371]), .A1N(n25410), .B0(n25395), .Y(n25396) );
  AOI22XL U16762 ( .A0(n3028), .A1(w1[275]), .B0(in_valid_w1), .B1(weight1[19]), .Y(n25395) );
  OAI2BB1XL U16763 ( .A0N(w1[372]), .A1N(n25410), .B0(n25387), .Y(n25388) );
  AOI22XL U16764 ( .A0(n3028), .A1(w1[276]), .B0(in_valid_w1), .B1(weight1[20]), .Y(n25387) );
  OAI2BB1XL U16765 ( .A0N(w1[373]), .A1N(n25410), .B0(n25374), .Y(n25375) );
  AOI22XL U16766 ( .A0(n3028), .A1(w1[277]), .B0(in_valid_w1), .B1(weight1[21]), .Y(n25374) );
  OAI2BB1XL U16767 ( .A0N(w1[375]), .A1N(n25410), .B0(n24323), .Y(n24324) );
  AOI22XL U16768 ( .A0(n3028), .A1(w1[279]), .B0(in_valid_w1), .B1(weight1[23]), .Y(n24323) );
  OAI2BB1XL U16769 ( .A0N(w1[376]), .A1N(n25410), .B0(n25121), .Y(n25122) );
  AOI22XL U16770 ( .A0(n3028), .A1(w1[280]), .B0(in_valid_w1), .B1(weight1[24]), .Y(n25121) );
  OAI2BB1XL U16771 ( .A0N(w1[377]), .A1N(n25410), .B0(n24368), .Y(n24369) );
  AOI22XL U16772 ( .A0(n3028), .A1(w1[281]), .B0(in_valid_w1), .B1(weight1[25]), .Y(n24368) );
  OAI2BB1XL U16773 ( .A0N(w1[378]), .A1N(n3052), .B0(n24061), .Y(n24062) );
  AOI22XL U16774 ( .A0(n3028), .A1(w1[282]), .B0(in_valid_w1), .B1(weight1[26]), .Y(n24061) );
  OAI2BB1XL U16775 ( .A0N(w1[381]), .A1N(n25410), .B0(n25111), .Y(n25112) );
  AOI22XL U16776 ( .A0(n3028), .A1(w1[285]), .B0(in_valid_w1), .B1(weight1[29]), .Y(n25111) );
  OAI2BB1XL U16777 ( .A0N(w1[382]), .A1N(n3052), .B0(n25843), .Y(n25844) );
  AOI22XL U16778 ( .A0(n3064), .A1(w1[286]), .B0(in_valid_w1), .B1(weight1[30]), .Y(n25843) );
  MXI2XL U16779 ( .A(data[0]), .B(data[32]), .S0(n3229), .Y(n1614) );
  MXI2XL U16780 ( .A(data[1]), .B(data[33]), .S0(n3229), .Y(n1615) );
  MXI2XL U16781 ( .A(data[2]), .B(data[34]), .S0(n3229), .Y(n1616) );
  MXI2XL U16782 ( .A(data[3]), .B(data[35]), .S0(n4579), .Y(n1617) );
  MXI2XL U16783 ( .A(data[4]), .B(data[36]), .S0(n4579), .Y(n1618) );
  MXI2XL U16784 ( .A(data[5]), .B(data[37]), .S0(n3123), .Y(n1619) );
  MXI2XL U16785 ( .A(data[6]), .B(data[38]), .S0(n3123), .Y(n1620) );
  MXI2XL U16786 ( .A(data[7]), .B(data[39]), .S0(n3123), .Y(n1621) );
  MXI2XL U16787 ( .A(data[8]), .B(data[40]), .S0(n4579), .Y(n1622) );
  MXI2XL U16788 ( .A(data[9]), .B(data[41]), .S0(n3229), .Y(n1623) );
  MXI2XL U16789 ( .A(data[10]), .B(data[42]), .S0(n3123), .Y(n1624) );
  MXI2XL U16790 ( .A(data[11]), .B(data[43]), .S0(n3229), .Y(n1625) );
  MXI2XL U16791 ( .A(data[12]), .B(data[44]), .S0(n3229), .Y(n1626) );
  MXI2XL U16792 ( .A(data[13]), .B(data[45]), .S0(n3123), .Y(n1627) );
  MXI2XL U16793 ( .A(data[14]), .B(data[46]), .S0(n3123), .Y(n1628) );
  MXI2XL U16794 ( .A(data[15]), .B(data[47]), .S0(n3229), .Y(n1629) );
  MXI2XL U16795 ( .A(data[16]), .B(data[48]), .S0(n3123), .Y(n1630) );
  MXI2XL U16796 ( .A(data[17]), .B(data[49]), .S0(n3229), .Y(n1631) );
  MXI2XL U16797 ( .A(data[18]), .B(data[50]), .S0(n3229), .Y(n1632) );
  MXI2XL U16798 ( .A(data[19]), .B(data[51]), .S0(n3229), .Y(n1633) );
  MXI2XL U16799 ( .A(data[20]), .B(data[52]), .S0(n3123), .Y(n1634) );
  MXI2XL U16800 ( .A(data[21]), .B(data[53]), .S0(n3229), .Y(n1635) );
  MXI2XL U16801 ( .A(data[22]), .B(data[54]), .S0(n4579), .Y(n1636) );
  MXI2XL U16802 ( .A(data[23]), .B(data[55]), .S0(n3123), .Y(n1637) );
  MXI2XL U16803 ( .A(data[25]), .B(data[57]), .S0(n3123), .Y(n1639) );
  MXI2XL U16804 ( .A(data[27]), .B(data[59]), .S0(n3123), .Y(n1641) );
  MXI2XL U16805 ( .A(data[29]), .B(data[61]), .S0(n3229), .Y(n1643) );
  MXI2XL U16806 ( .A(data[31]), .B(data[63]), .S0(n3123), .Y(n1645) );
  MXI2XL U16807 ( .A(data[55]), .B(data[87]), .S0(n3229), .Y(n1669) );
  MXI2XL U16808 ( .A(data[56]), .B(data[88]), .S0(n4579), .Y(n1670) );
  MXI2XL U16809 ( .A(data[57]), .B(data[89]), .S0(n4579), .Y(n1671) );
  MXI2XL U16810 ( .A(data[59]), .B(data[91]), .S0(n4579), .Y(n1673) );
  MXI2XL U16811 ( .A(data[60]), .B(data[92]), .S0(n4579), .Y(n1674) );
  MXI2XL U16812 ( .A(data[61]), .B(data[93]), .S0(n4579), .Y(n1675) );
  MXI2XL U16813 ( .A(data[63]), .B(data[95]), .S0(n3229), .Y(n1677) );
  MXI2XL U16814 ( .A(data[89]), .B(data[121]), .S0(n3123), .Y(n1703) );
  MXI2XL U16815 ( .A(data[91]), .B(data[123]), .S0(in_valid_d), .Y(n1705) );
  MXI2XL U16816 ( .A(data[92]), .B(data[124]), .S0(n3123), .Y(n1706) );
  MXI2XL U16817 ( .A(data[93]), .B(data[125]), .S0(n4579), .Y(n1707) );
  MXI2XL U16818 ( .A(data[95]), .B(data[127]), .S0(n4579), .Y(n1709) );
  INVXL U16819 ( .A(n24022), .Y(n24023) );
  INVXL U16820 ( .A(n25216), .Y(n25217) );
  INVXL U16821 ( .A(n25213), .Y(n25214) );
  INVXL U16822 ( .A(n25210), .Y(n25211) );
  MXI2XL U16823 ( .A(data[127]), .B(data_point[31]), .S0(n4579), .Y(n1741) );
  OAI211XL U16824 ( .A0(iter[2]), .A1(n23062), .B0(n23985), .C0(n23055), .Y(
        n1743) );
  OAI211XL U16825 ( .A0(iter[4]), .A1(n23054), .B0(n23985), .C0(n23058), .Y(
        n1745) );
  OAI211XL U16826 ( .A0(iter[6]), .A1(n23057), .B0(n23985), .C0(n23060), .Y(
        n1747) );
  AOI222XL U16827 ( .A0(n23088), .A1(w1[65]), .B0(n3023), .B1(w1[33]), .C0(
        w1[161]), .C1(n3216), .Y(n1756) );
  AOI222XL U16828 ( .A0(n25567), .A1(w1[98]), .B0(n3023), .B1(w1[66]), .C0(
        w1[194]), .C1(n3216), .Y(n1761) );
  AOI222XL U16829 ( .A0(n23088), .A1(w1[99]), .B0(n3023), .B1(w1[67]), .C0(
        w1[195]), .C1(n3216), .Y(n1765) );
  AOI222XL U16830 ( .A0(n25567), .A1(w1[68]), .B0(n3023), .B1(w1[36]), .C0(
        w1[164]), .C1(n3216), .Y(n1768) );
  AOI222XL U16831 ( .A0(n23088), .A1(w1[36]), .B0(n3023), .B1(w1[4]), .C0(
        w1[132]), .C1(n3216), .Y(n1771) );
  AOI222XL U16832 ( .A0(n23088), .A1(w1[70]), .B0(n3023), .B1(w1[38]), .C0(
        w1[166]), .C1(n3216), .Y(n1776) );
  AOI222XL U16833 ( .A0(n25567), .A1(w1[38]), .B0(n3023), .B1(w1[6]), .C0(
        w1[134]), .C1(n3216), .Y(n1779) );
  AOI222XL U16834 ( .A0(n23088), .A1(w1[71]), .B0(n3023), .B1(w1[39]), .C0(
        w1[167]), .C1(n3216), .Y(n1780) );
  AOI222XL U16835 ( .A0(n3061), .A1(w1[103]), .B0(n3023), .B1(w1[71]), .C0(
        w1[199]), .C1(n3216), .Y(n1781) );
  AOI222XL U16836 ( .A0(n25567), .A1(w1[39]), .B0(n3023), .B1(w1[7]), .C0(
        w1[135]), .C1(n3216), .Y(n1783) );
  AOI222XL U16837 ( .A0(n23088), .A1(w1[72]), .B0(n3023), .B1(w1[40]), .C0(
        w1[168]), .C1(n3216), .Y(n1784) );
  AOI222XL U16838 ( .A0(n25567), .A1(w1[104]), .B0(n3023), .B1(w1[72]), .C0(
        w1[200]), .C1(n3216), .Y(n1785) );
  AOI222XL U16839 ( .A0(n23088), .A1(w1[40]), .B0(n3023), .B1(w1[8]), .C0(
        w1[136]), .C1(n3216), .Y(n1787) );
  AOI222XL U16840 ( .A0(n25567), .A1(w1[73]), .B0(n3023), .B1(w1[41]), .C0(
        w1[169]), .C1(n3216), .Y(n1788) );
  AOI222XL U16841 ( .A0(n25567), .A1(w1[105]), .B0(n3023), .B1(w1[73]), .C0(
        w1[201]), .C1(n3216), .Y(n1789) );
  AOI222XL U16842 ( .A0(n3061), .A1(w1[42]), .B0(n3023), .B1(w1[10]), .C0(
        w1[138]), .C1(n3216), .Y(n1795) );
  AOI222XL U16843 ( .A0(n23088), .A1(w1[75]), .B0(n3051), .B1(w1[43]), .C0(
        w1[171]), .C1(n3216), .Y(n1796) );
  AOI222XL U16844 ( .A0(n23088), .A1(w1[107]), .B0(n3051), .B1(w1[75]), .C0(
        w1[203]), .C1(n3216), .Y(n1797) );
  AOI222XL U16845 ( .A0(n25567), .A1(w1[43]), .B0(n3051), .B1(w1[11]), .C0(
        w1[139]), .C1(n3216), .Y(n1799) );
  AOI222XL U16846 ( .A0(n25567), .A1(w1[77]), .B0(n3051), .B1(w1[45]), .C0(
        w1[173]), .C1(n3216), .Y(n1804) );
  AOI222XL U16847 ( .A0(n25567), .A1(w1[109]), .B0(n3051), .B1(w1[77]), .C0(
        w1[205]), .C1(n3216), .Y(n1805) );
  AOI222XL U16848 ( .A0(n23088), .A1(w1[45]), .B0(n3051), .B1(w1[13]), .C0(
        w1[141]), .C1(n3216), .Y(n1807) );
  AOI222XL U16849 ( .A0(n25567), .A1(w1[110]), .B0(n3051), .B1(w1[78]), .C0(
        w1[206]), .C1(n3216), .Y(n1809) );
  AOI222XL U16850 ( .A0(n23088), .A1(w1[79]), .B0(n3051), .B1(w1[47]), .C0(
        w1[175]), .C1(n3216), .Y(n1812) );
  AOI222XL U16851 ( .A0(n3061), .A1(w1[111]), .B0(n3051), .B1(w1[79]), .C0(
        w1[207]), .C1(n3216), .Y(n1813) );
  AOI222XL U16852 ( .A0(n25567), .A1(w1[47]), .B0(n3051), .B1(w1[15]), .C0(
        w1[143]), .C1(n3216), .Y(n1815) );
  AOI222XL U16853 ( .A0(n25567), .A1(w1[48]), .B0(n3051), .B1(w1[16]), .C0(
        w1[144]), .C1(n3216), .Y(n1819) );
  AOI222XL U16854 ( .A0(n23088), .A1(w1[113]), .B0(n3051), .B1(w1[81]), .C0(
        w1[209]), .C1(n3216), .Y(n1821) );
  AOI222XL U16855 ( .A0(n25567), .A1(w1[82]), .B0(n3051), .B1(w1[50]), .C0(
        w1[178]), .C1(n3216), .Y(n1824) );
  AOI222XL U16856 ( .A0(n25567), .A1(w1[50]), .B0(n3051), .B1(w1[18]), .C0(
        w1[146]), .C1(n3216), .Y(n1827) );
  AOI222XL U16857 ( .A0(n25567), .A1(w1[51]), .B0(n3051), .B1(w1[19]), .C0(
        w1[147]), .C1(n3216), .Y(n1831) );
  AOI222XL U16858 ( .A0(n23088), .A1(w1[84]), .B0(n3051), .B1(w1[52]), .C0(
        w1[180]), .C1(n3216), .Y(n1832) );
  AOI222XL U16859 ( .A0(n25567), .A1(w1[116]), .B0(n3051), .B1(w1[84]), .C0(
        w1[212]), .C1(n3216), .Y(n1833) );
  AOI222XL U16860 ( .A0(n25567), .A1(w1[52]), .B0(n3051), .B1(w1[20]), .C0(
        w1[148]), .C1(n3216), .Y(n1835) );
  AOI222XL U16861 ( .A0(n25567), .A1(w1[85]), .B0(n3051), .B1(w1[53]), .C0(
        w1[181]), .C1(n3216), .Y(n1836) );
  AOI222XL U16862 ( .A0(n25567), .A1(w1[117]), .B0(n3051), .B1(w1[85]), .C0(
        w1[213]), .C1(n3216), .Y(n1837) );
  AOI222XL U16863 ( .A0(n25567), .A1(w1[53]), .B0(n3051), .B1(w1[21]), .C0(
        w1[149]), .C1(n3216), .Y(n1839) );
  AOI222XL U16864 ( .A0(n25567), .A1(w1[86]), .B0(n3051), .B1(w1[54]), .C0(
        w1[182]), .C1(n25541), .Y(n1840) );
  AOI222XL U16865 ( .A0(n23088), .A1(w1[54]), .B0(n3051), .B1(w1[22]), .C0(
        w1[150]), .C1(n3216), .Y(n1843) );
  AOI222XL U16866 ( .A0(n25567), .A1(w1[87]), .B0(n3216), .B1(w1[183]), .C0(
        w1[55]), .C1(n25410), .Y(n1844) );
  AOI222XL U16867 ( .A0(n23088), .A1(w1[119]), .B0(n3216), .B1(w1[215]), .C0(
        w1[87]), .C1(n25410), .Y(n1845) );
  AOI222XL U16868 ( .A0(n25567), .A1(w1[55]), .B0(w1[23]), .B1(n3052), .C0(
        w1[151]), .C1(n3216), .Y(n1847) );
  AOI222XL U16869 ( .A0(n25567), .A1(w1[88]), .B0(n3216), .B1(w1[184]), .C0(
        w1[56]), .C1(n25410), .Y(n1848) );
  AOI222XL U16870 ( .A0(n25567), .A1(w1[120]), .B0(n3216), .B1(w1[216]), .C0(
        w1[88]), .C1(n25410), .Y(n1849) );
  AOI222XL U16871 ( .A0(n23088), .A1(w1[56]), .B0(w1[24]), .B1(n25410), .C0(
        w1[152]), .C1(n3216), .Y(n1851) );
  AOI222XL U16872 ( .A0(n25567), .A1(w1[89]), .B0(n3216), .B1(w1[185]), .C0(
        w1[57]), .C1(n25410), .Y(n1852) );
  AOI222XL U16873 ( .A0(n25567), .A1(w1[121]), .B0(n3216), .B1(w1[217]), .C0(
        w1[89]), .C1(n25410), .Y(n1853) );
  AOI222XL U16874 ( .A0(n3061), .A1(w1[57]), .B0(w1[25]), .B1(n4576), .C0(
        w1[153]), .C1(n3216), .Y(n1855) );
  AOI222XL U16875 ( .A0(n3061), .A1(w1[90]), .B0(n3216), .B1(w1[186]), .C0(
        w1[58]), .C1(n25410), .Y(n1856) );
  AOI222XL U16876 ( .A0(n3061), .A1(w1[122]), .B0(n3216), .B1(w1[218]), .C0(
        w1[90]), .C1(n3023), .Y(n1857) );
  AOI222XL U16877 ( .A0(n3061), .A1(w1[58]), .B0(w1[26]), .B1(n25410), .C0(
        w1[154]), .C1(n3216), .Y(n1859) );
  AOI222XL U16878 ( .A0(n23088), .A1(w1[123]), .B0(n3216), .B1(w1[219]), .C0(
        w1[91]), .C1(n25410), .Y(n1861) );
  AOI222XL U16879 ( .A0(n3061), .A1(w1[92]), .B0(n3216), .B1(w1[188]), .C0(
        w1[60]), .C1(n25410), .Y(n1864) );
  AOI222XL U16880 ( .A0(n3061), .A1(w1[124]), .B0(n3216), .B1(w1[220]), .C0(
        w1[92]), .C1(n25410), .Y(n1865) );
  AOI222XL U16881 ( .A0(n23088), .A1(w1[60]), .B0(w1[28]), .B1(n4576), .C0(
        w1[156]), .C1(n3216), .Y(n1867) );
  AOI222XL U16882 ( .A0(n3061), .A1(w1[125]), .B0(n3216), .B1(w1[221]), .C0(
        w1[93]), .C1(n25410), .Y(n1869) );
  AOI222XL U16883 ( .A0(n3061), .A1(w1[94]), .B0(n3216), .B1(w1[190]), .C0(
        w1[62]), .C1(n25410), .Y(n1872) );
  AOI222XL U16884 ( .A0(n3061), .A1(w1[126]), .B0(n3216), .B1(w1[222]), .C0(
        w1[94]), .C1(n25410), .Y(n1873) );
  AOI222XL U16885 ( .A0(n3061), .A1(w1[62]), .B0(w1[30]), .B1(n4576), .C0(
        w1[158]), .C1(n3216), .Y(n1875) );
  AOI222XL U16886 ( .A0(n23088), .A1(w1[95]), .B0(n3216), .B1(w1[191]), .C0(
        w1[63]), .C1(n25410), .Y(n1876) );
  AOI222XL U16887 ( .A0(n3061), .A1(w1[127]), .B0(n3216), .B1(w1[223]), .C0(
        w1[95]), .C1(n25410), .Y(n1877) );
  AOI222XL U16888 ( .A0(n3061), .A1(w1[63]), .B0(n3216), .B1(w1[159]), .C0(
        n3052), .C1(w1[31]), .Y(n1879) );
  AOI222XL U16889 ( .A0(n23088), .A1(w1[160]), .B0(n3051), .B1(w1[128]), .C0(
        w1[256]), .C1(n3216), .Y(n1883) );
  AOI222XL U16890 ( .A0(n3061), .A1(w1[193]), .B0(n3051), .B1(w1[161]), .C0(
        w1[289]), .C1(n3216), .Y(n1884) );
  AOI222XL U16891 ( .A0(n3061), .A1(w1[161]), .B0(n3051), .B1(w1[129]), .C0(
        w1[257]), .C1(n3216), .Y(n1887) );
  AOI222XL U16892 ( .A0(n3061), .A1(w1[162]), .B0(n3051), .B1(w1[130]), .C0(
        w1[258]), .C1(n3216), .Y(n1891) );
  AOI222XL U16893 ( .A0(n3061), .A1(w1[195]), .B0(n3051), .B1(w1[163]), .C0(
        w1[291]), .C1(n3216), .Y(n1892) );
  AOI222XL U16894 ( .A0(n3061), .A1(w1[163]), .B0(n3051), .B1(w1[131]), .C0(
        w1[259]), .C1(n3216), .Y(n1895) );
  AOI222XL U16895 ( .A0(n3061), .A1(w1[196]), .B0(n3113), .B1(w1[164]), .C0(
        w1[292]), .C1(n3216), .Y(n1896) );
  AOI222XL U16896 ( .A0(n3061), .A1(w1[164]), .B0(n3113), .B1(w1[132]), .C0(
        w1[260]), .C1(n3216), .Y(n1899) );
  AOI222XL U16897 ( .A0(n3061), .A1(w1[197]), .B0(n3113), .B1(w1[165]), .C0(
        w1[293]), .C1(n3216), .Y(n1900) );
  AOI222XL U16898 ( .A0(n3061), .A1(w1[165]), .B0(n3113), .B1(w1[133]), .C0(
        w1[261]), .C1(n3216), .Y(n1903) );
  AOI222XL U16899 ( .A0(n3061), .A1(w1[198]), .B0(n3113), .B1(w1[166]), .C0(
        w1[294]), .C1(n3216), .Y(n1904) );
  AOI222XL U16900 ( .A0(n3061), .A1(w1[166]), .B0(n3113), .B1(w1[134]), .C0(
        w1[262]), .C1(n3216), .Y(n1907) );
  AOI222XL U16901 ( .A0(n3061), .A1(w1[199]), .B0(n3113), .B1(w1[167]), .C0(
        w1[295]), .C1(n3216), .Y(n1908) );
  AOI222XL U16902 ( .A0(n23088), .A1(w1[167]), .B0(n3113), .B1(w1[135]), .C0(
        w1[263]), .C1(n3216), .Y(n1911) );
  AOI222XL U16903 ( .A0(n23088), .A1(w1[203]), .B0(n3113), .B1(w1[171]), .C0(
        w1[299]), .C1(n3216), .Y(n1924) );
  AOI222XL U16904 ( .A0(n3061), .A1(w1[171]), .B0(n3113), .B1(w1[139]), .C0(
        w1[267]), .C1(n3216), .Y(n1927) );
  AOI222XL U16905 ( .A0(n3061), .A1(w1[172]), .B0(n3113), .B1(w1[140]), .C0(
        w1[268]), .C1(n3216), .Y(n1931) );
  AOI222XL U16906 ( .A0(n3061), .A1(w1[173]), .B0(n3113), .B1(w1[141]), .C0(
        w1[269]), .C1(n3216), .Y(n1935) );
  AOI222XL U16907 ( .A0(n3061), .A1(w1[206]), .B0(n3113), .B1(w1[174]), .C0(
        w1[302]), .C1(n3216), .Y(n1936) );
  AOI222XL U16908 ( .A0(n3061), .A1(w1[174]), .B0(n3113), .B1(w1[142]), .C0(
        w1[270]), .C1(n3216), .Y(n1939) );
  AOI222XL U16909 ( .A0(n3061), .A1(w1[207]), .B0(n3113), .B1(w1[175]), .C0(
        w1[303]), .C1(n3216), .Y(n1940) );
  AOI222XL U16910 ( .A0(n3061), .A1(w1[175]), .B0(n3113), .B1(w1[143]), .C0(
        w1[271]), .C1(n3216), .Y(n1943) );
  AOI222XL U16911 ( .A0(n3061), .A1(w1[240]), .B0(n3113), .B1(w1[208]), .C0(
        w1[336]), .C1(n3216), .Y(n1945) );
  AOI222XL U16912 ( .A0(n23088), .A1(w1[209]), .B0(n3113), .B1(w1[177]), .C0(
        w1[305]), .C1(n3216), .Y(n1948) );
  AOI222XL U16913 ( .A0(n3061), .A1(w1[177]), .B0(n3113), .B1(w1[145]), .C0(
        w1[273]), .C1(n3216), .Y(n1951) );
  AOI222XL U16914 ( .A0(n3061), .A1(w1[178]), .B0(n3113), .B1(w1[146]), .C0(
        w1[274]), .C1(n3216), .Y(n1955) );
  AOI222XL U16915 ( .A0(n23088), .A1(w1[212]), .B0(n3113), .B1(w1[180]), .C0(
        w1[308]), .C1(n3216), .Y(n1960) );
  AOI222XL U16916 ( .A0(n3061), .A1(w1[180]), .B0(n3113), .B1(w1[148]), .C0(
        w1[276]), .C1(n3216), .Y(n1963) );
  AOI222XL U16917 ( .A0(n3061), .A1(w1[213]), .B0(n4578), .B1(w1[181]), .C0(
        w1[309]), .C1(n3216), .Y(n1964) );
  AOI222XL U16918 ( .A0(n3061), .A1(w1[181]), .B0(n3051), .B1(w1[149]), .C0(
        w1[277]), .C1(n3216), .Y(n1967) );
  AOI222XL U16919 ( .A0(n3061), .A1(w1[214]), .B0(n3051), .B1(w1[182]), .C0(
        w1[310]), .C1(n3216), .Y(n1968) );
  AOI222XL U16920 ( .A0(n3061), .A1(w1[182]), .B0(n3051), .B1(w1[150]), .C0(
        w1[278]), .C1(n3216), .Y(n1971) );
  AOI222XL U16921 ( .A0(n3061), .A1(w1[215]), .B0(n3051), .B1(w1[183]), .C0(
        w1[311]), .C1(n3216), .Y(n1972) );
  AOI222XL U16922 ( .A0(n3061), .A1(w1[183]), .B0(w1[279]), .B1(n3216), .C0(
        w1[151]), .C1(n25410), .Y(n1975) );
  AOI222XL U16923 ( .A0(n3061), .A1(w1[216]), .B0(n3023), .B1(w1[184]), .C0(
        w1[312]), .C1(n3216), .Y(n1976) );
  AOI222XL U16924 ( .A0(n3061), .A1(w1[184]), .B0(w1[280]), .B1(n3216), .C0(
        w1[152]), .C1(n25410), .Y(n1979) );
  AOI222XL U16925 ( .A0(n3061), .A1(w1[185]), .B0(w1[281]), .B1(n3216), .C0(
        w1[153]), .C1(n25410), .Y(n1983) );
  AOI222XL U16926 ( .A0(n3061), .A1(w1[186]), .B0(w1[282]), .B1(n3216), .C0(
        w1[154]), .C1(n25410), .Y(n1987) );
  AOI222XL U16927 ( .A0(n3061), .A1(w1[187]), .B0(w1[283]), .B1(n3216), .C0(
        w1[155]), .C1(n25410), .Y(n1991) );
  AOI222XL U16928 ( .A0(n23088), .A1(w1[220]), .B0(n3051), .B1(w1[188]), .C0(
        w1[316]), .C1(n3216), .Y(n1992) );
  AOI222XL U16929 ( .A0(n3061), .A1(w1[188]), .B0(w1[284]), .B1(n3216), .C0(
        w1[156]), .C1(n25410), .Y(n1995) );
  AOI222XL U16930 ( .A0(n3061), .A1(w1[221]), .B0(n3051), .B1(w1[189]), .C0(
        w1[317]), .C1(n3216), .Y(n1996) );
  AOI222XL U16931 ( .A0(n3061), .A1(w1[189]), .B0(w1[285]), .B1(n3216), .C0(
        w1[157]), .C1(n25410), .Y(n1999) );
  AOI222XL U16932 ( .A0(n3061), .A1(w1[190]), .B0(w1[286]), .B1(n3216), .C0(
        w1[158]), .C1(n25410), .Y(n2003) );
  AOI222XL U16933 ( .A0(n3061), .A1(w1[223]), .B0(n3051), .B1(w1[191]), .C0(
        w1[319]), .C1(n3216), .Y(n2004) );
  INVXL U16934 ( .A(n23355), .Y(n23356) );
  INVXL U16935 ( .A(n23324), .Y(n23325) );
  OAI31XL U16936 ( .A0(n22468), .A1(n3226), .A2(n23235), .B0(n22467), .Y(
        n22469) );
  AOI22XL U16937 ( .A0(n3052), .A1(w1[278]), .B0(w1[310]), .B1(n3061), .Y(
        n22467) );
  INVXL U16938 ( .A(n23041), .Y(n22468) );
  AOI222XL U16939 ( .A0(n3061), .A1(w1[319]), .B0(n3216), .B1(n23137), .C0(
        w1[287]), .C1(n25410), .Y(n2135) );
  AOI222XL U16940 ( .A0(n25659), .A1(n25292), .B0(w2[95]), .B1(n25822), .C0(
        in_valid_w2), .C1(weight2[31]), .Y(n2231) );
  AOI21XL U16941 ( .A0(n23355), .A1(n23429), .B0(n23259), .Y(n23260) );
  OAI22XL U16942 ( .A0(n23039), .A1(target_temp[0]), .B0(target[0]), .B1(
        n17167), .Y(n23259) );
  INVXL U16943 ( .A(n23254), .Y(n2236) );
  OAI22XL U16944 ( .A0(n23039), .A1(target_temp[4]), .B0(target[4]), .B1(
        n15940), .Y(n23253) );
  AOI222XL U16945 ( .A0(n23234), .A1(n23429), .B0(target_temp[27]), .B1(n23428), .C0(in_valid_t), .C1(target[27]), .Y(n2259) );
  OAI31XL U16946 ( .A0(learning_rate[23]), .A1(n23985), .A2(n22471), .B0(
        n22470), .Y(n2628) );
  NAND3XL U16947 ( .A(n24015), .B(n24008), .C(n24004), .Y(n24005) );
  AOI2BB1XL U16948 ( .A0N(n21102), .A1N(n22471), .B0(n24007), .Y(n21103) );
  OAI22XL U16949 ( .A0(n25856), .A1(n23053), .B0(n23052), .B1(n23982), .Y(
        n2624) );
  AOI21XL U16950 ( .A0(n24009), .A1(n24008), .B0(n24007), .Y(n24010) );
  INVXL U16951 ( .A(n23643), .Y(n23636) );
  XOR2XL U16952 ( .A(n25133), .B(n25136), .Y(n25134) );
  NOR3XL U16953 ( .A(n25258), .B(n25257), .C(n3121), .Y(n25259) );
  OAI21XL U16954 ( .A0(n24315), .A1(n3121), .B0(n5355), .Y(n2570) );
  AOI21XL U16955 ( .A0(n23972), .A1(in_valid_d), .B0(n5356), .Y(n5355) );
  AOI22XL U16956 ( .A0(n23717), .A1(n3223), .B0(n25723), .B1(temp0[23]), .Y(
        n23719) );
  OAI211XL U16957 ( .A0(n25829), .A1(n23680), .B0(n25699), .C0(n23679), .Y(
        n23681) );
  AOI211XL U16958 ( .A0(n25691), .A1(in_valid_d), .B0(n25248), .C0(n25247), 
        .Y(n25249) );
  AOI211XL U16959 ( .A0(n25245), .A1(n25244), .B0(n3115), .C0(n25242), .Y(
        n25248) );
  NOR2XL U16960 ( .A(n25837), .B(n25246), .Y(n25247) );
  AOI22XL U16961 ( .A0(n25668), .A1(n25667), .B0(n2982), .B1(temp1[31]), .Y(
        n25669) );
  NOR2XL U16962 ( .A(n25666), .B(n3121), .Y(n25667) );
  BUFX3 U16963 ( .A(n11479), .Y(n5770) );
  BUFX3 U16964 ( .A(n11479), .Y(n4875) );
  INVX4 U16965 ( .A(n4622), .Y(n19542) );
  XOR2X1 U16966 ( .A(n5391), .B(M1_b_15_), .Y(n6208) );
  CLKINVX3 U16967 ( .A(n13791), .Y(n13045) );
  XNOR2X1 U16968 ( .A(n19382), .B(n19381), .Y(n4622) );
  NAND2X4 U16969 ( .A(n3046), .B(n6292), .Y(n4592) );
  NAND2X1 U16970 ( .A(n17350), .B(n17349), .Y(n4595) );
  NAND2X1 U16971 ( .A(n17344), .B(n17342), .Y(n4598) );
  CLKINVX3 U16972 ( .A(M3_mult_x_15_b_20_), .Y(n6112) );
  AOI2BB1X2 U16973 ( .A0N(n7382), .A1N(n26008), .B0(n5566), .Y(n6476) );
  NOR2X2 U16974 ( .A(n4583), .B(n6224), .Y(n25149) );
  AND2X2 U16975 ( .A(n10736), .B(n4673), .Y(n4599) );
  INVX4 U16976 ( .A(n7615), .Y(n23221) );
  INVX1 U16977 ( .A(n25813), .Y(n5434) );
  INVX1 U16978 ( .A(n24293), .Y(n4790) );
  AND2X1 U16979 ( .A(n10215), .B(n10214), .Y(n4602) );
  AND2X1 U16980 ( .A(n10239), .B(n10238), .Y(n4606) );
  XOR2X1 U16981 ( .A(n23409), .B(n21455), .Y(n21507) );
  BUFX3 U16982 ( .A(M2_b_16_), .Y(n10335) );
  NOR2X2 U16983 ( .A(n18890), .B(n18886), .Y(n18865) );
  XOR2X2 U16984 ( .A(n21454), .B(n21453), .Y(n21580) );
  XNOR2X2 U16985 ( .A(n4785), .B(M5_a_8_), .Y(n16943) );
  BUFX3 U16986 ( .A(n16943), .Y(n16688) );
  INVX1 U16987 ( .A(n12387), .Y(n4961) );
  CLKINVX3 U16988 ( .A(n5583), .Y(n7146) );
  OR2X2 U16989 ( .A(n10472), .B(n10471), .Y(n4619) );
  OR2X2 U16990 ( .A(n18307), .B(n18306), .Y(n4620) );
  CLKBUFX8 U16991 ( .A(n11496), .Y(M3_mult_x_15_b_1_) );
  CLKINVX3 U16992 ( .A(n14081), .Y(n13173) );
  BUFX3 U16993 ( .A(n6223), .Y(n5604) );
  XNOR2X1 U16994 ( .A(n14973), .B(n14972), .Y(n15161) );
  AND2X2 U16995 ( .A(n10321), .B(n10463), .Y(n4626) );
  BUFX3 U16996 ( .A(n13898), .Y(n4848) );
  NAND2X1 U16997 ( .A(n17339), .B(n17338), .Y(n4632) );
  CLKBUFX8 U16998 ( .A(M3_mult_x_15_b_14_), .Y(n12701) );
  AND2X1 U16999 ( .A(n13465), .B(n13464), .Y(n4633) );
  OR2X2 U17000 ( .A(n17130), .B(n17129), .Y(n4634) );
  CLKBUFX8 U17001 ( .A(n11628), .Y(n12718) );
  NAND2X2 U17002 ( .A(n11529), .B(n9080), .Y(n10337) );
  INVX1 U17003 ( .A(n10337), .Y(n6140) );
  OAI21X1 U17004 ( .A0(n25813), .A1(n26266), .B0(n17479), .Y(M4_a_0_) );
  OR2X2 U17005 ( .A(n6662), .B(n6661), .Y(n4635) );
  INVX1 U17006 ( .A(n17225), .Y(n17303) );
  XNOR2X1 U17007 ( .A(M4_a_20_), .B(M4_a_19_), .Y(n17605) );
  CLKINVX3 U17008 ( .A(n25269), .Y(n15764) );
  NAND2X4 U17009 ( .A(n6289), .B(n6745), .Y(n4642) );
  NOR2X1 U17010 ( .A(n17107), .B(n17106), .Y(n17315) );
  INVX1 U17011 ( .A(n10503), .Y(n10619) );
  OR2X2 U17012 ( .A(n14080), .B(n13169), .Y(n4644) );
  AND4X2 U17013 ( .A(n24066), .B(n20173), .C(n20194), .D(n20172), .Y(n24692)
         );
  OR2X2 U17014 ( .A(n12985), .B(n12991), .Y(n4647) );
  XOR2X1 U17015 ( .A(M3_mult_x_15_n1682), .B(n18428), .Y(n4649) );
  INVX1 U17016 ( .A(n18928), .Y(n18938) );
  INVX1 U17017 ( .A(n13025), .Y(n17457) );
  AND2X2 U17018 ( .A(n5899), .B(n19044), .Y(n4651) );
  CLKINVX3 U17019 ( .A(n5033), .Y(n20700) );
  INVX1 U17020 ( .A(M3_mult_x_15_b_1_), .Y(n5705) );
  NOR2X1 U17021 ( .A(n13984), .B(n13983), .Y(n14637) );
  INVX1 U17022 ( .A(n20312), .Y(n4944) );
  OR3XL U17023 ( .A(n12940), .B(n24040), .C(n11622), .Y(n4656) );
  AND2X2 U17024 ( .A(n17908), .B(n4882), .Y(n17919) );
  XNOR3X2 U17025 ( .A(n4990), .B(n11891), .C(n11890), .Y(n4658) );
  CLKINVX3 U17026 ( .A(n5667), .Y(n17375) );
  OR2X2 U17027 ( .A(n6274), .B(n25993), .Y(n4662) );
  XNOR2X1 U17028 ( .A(n11972), .B(n11973), .Y(n4666) );
  XNOR2X1 U17029 ( .A(n14156), .B(n5488), .Y(n4667) );
  INVX1 U17030 ( .A(n12689), .Y(n6114) );
  ADDFX2 U17031 ( .A(n12656), .B(n12655), .CI(n12654), .CO(n12689), .S(n12678)
         );
  AND2X2 U17032 ( .A(n20671), .B(n20670), .Y(n4671) );
  OR2X2 U17033 ( .A(n11483), .B(n6166), .Y(n4674) );
  CLKINVX3 U17034 ( .A(M2_a_5_), .Y(n9878) );
  INVX4 U17035 ( .A(n7534), .Y(n23220) );
  NAND2X2 U17036 ( .A(n13039), .B(n5158), .Y(n23174) );
  OR2XL U17037 ( .A(M3_mult_x_15_a_17_), .B(n4945), .Y(n4693) );
  INVX4 U17038 ( .A(n7711), .Y(n23219) );
  OR2XL U17039 ( .A(n5677), .B(n17039), .Y(n4694) );
  NAND2X1 U17040 ( .A(n12823), .B(n12822), .Y(n4695) );
  NOR2X1 U17041 ( .A(n20654), .B(n20653), .Y(n4698) );
  CLKINVX3 U17042 ( .A(n3202), .Y(n5957) );
  AND2X1 U17043 ( .A(n23997), .B(n3027), .Y(n4710) );
  OR2XL U17044 ( .A(n23884), .B(n26529), .Y(n4711) );
  CLKINVX2 U17045 ( .A(n3227), .Y(n25696) );
  XNOR2X1 U17046 ( .A(n15970), .B(n16884), .Y(n16684) );
  XOR2X2 U17047 ( .A(n20924), .B(n20923), .Y(n20933) );
  BUFX3 U17048 ( .A(n11482), .Y(M3_mult_x_15_b_22_) );
  XOR2X2 U17049 ( .A(n19014), .B(n18864), .Y(n18972) );
  OAI22XL U17050 ( .A0(n7535), .A1(n7038), .B0(n7049), .B1(n7460), .Y(n7043)
         );
  AOI22X2 U17051 ( .A0(n19079), .A1(n3139), .B0(n3455), .B1(n20956), .Y(n23770) );
  ADDFHX1 U17052 ( .A(n9244), .B(n9243), .CI(n9242), .CO(n9290), .S(n9256) );
  ADDFHX1 U17053 ( .A(n9375), .B(n9374), .CI(n9373), .CO(n9328), .S(n9412) );
  NAND2X2 U17054 ( .A(n13988), .B(n13987), .Y(n14632) );
  CLKINVX3 U17055 ( .A(n14119), .Y(n14156) );
  XOR2X1 U17056 ( .A(n14196), .B(n5512), .Y(n13698) );
  OAI21X1 U17057 ( .A0(n25747), .A1(n3024), .B0(n25746), .Y(n25748) );
  AOI22XL U17058 ( .A0(n19667), .A1(n19642), .B0(n19651), .B1(n19641), .Y(
        n19647) );
  AOI21XL U17059 ( .A0(n19729), .A1(n3036), .B0(n2996), .Y(n19667) );
  XNOR2X1 U17060 ( .A(n3047), .B(M3_mult_x_15_b_9_), .Y(n16540) );
  XNOR2X1 U17061 ( .A(n3047), .B(n3201), .Y(n16380) );
  XNOR2X1 U17062 ( .A(n3047), .B(n3202), .Y(n15956) );
  XNOR2XL U17063 ( .A(n3047), .B(M3_mult_x_15_b_13_), .Y(n16408) );
  OAI22X1 U17064 ( .A0(n6214), .A1(n4860), .B0(n25906), .B1(n25796), .Y(n11488) );
  AOI21XL U17065 ( .A0(n25220), .A1(n25222), .B0(n25219), .Y(n25221) );
  AOI21XL U17066 ( .A0(M2_a_22_), .A1(n10540), .B0(n5255), .Y(
        M2_U3_U1_enc_tree_0__1__10_) );
  XNOR2X4 U17067 ( .A(M2_a_22_), .B(n5298), .Y(n10659) );
  INVX1 U17068 ( .A(n25687), .Y(n25745) );
  NAND2X1 U17069 ( .A(n5395), .B(n4599), .Y(n5364) );
  OAI21XL U17070 ( .A0(n3605), .A1(n7706), .B0(n7705), .Y(n7720) );
  OAI21XL U17071 ( .A0(n3605), .A1(n7810), .B0(n7809), .Y(n7813) );
  NAND2X1 U17072 ( .A(n7437), .B(n5622), .Y(n5621) );
  NAND2X2 U17073 ( .A(n10240), .B(n10135), .Y(n10179) );
  XOR2X1 U17074 ( .A(n5255), .B(n5298), .Y(n5078) );
  INVX1 U17075 ( .A(n10190), .Y(n10228) );
  NAND2X1 U17076 ( .A(n3895), .B(n20969), .Y(n20971) );
  NAND3X1 U17077 ( .A(n24179), .B(n4220), .C(n25796), .Y(n5267) );
  OAI21XL U17078 ( .A0(n15655), .A1(n15648), .B0(n15652), .Y(n15651) );
  NOR2X2 U17079 ( .A(n23966), .B(n14979), .Y(n14977) );
  NOR2X1 U17080 ( .A(n15916), .B(n15638), .Y(n25138) );
  NAND2X4 U17081 ( .A(n10659), .B(n9221), .Y(n10660) );
  OAI22X1 U17082 ( .A0(n16942), .A1(n15979), .B0(n16943), .B1(n16020), .Y(
        n16025) );
  OAI222X2 U17083 ( .A0(n6180), .A1(n15941), .B0(n25897), .B1(n25796), .C0(
        n17167), .C1(n23995), .Y(n11489) );
  OAI222X4 U17084 ( .A0(n6196), .A1(n11483), .B0(n25903), .B1(n21167), .C0(
        n23998), .C1(n17167), .Y(n11499) );
  CLKINVX3 U17085 ( .A(n25693), .Y(n24525) );
  OAI22X1 U17086 ( .A0(n18522), .A1(n17509), .B0(n3195), .B1(n17508), .Y(
        n17565) );
  XOR2X1 U17087 ( .A(n11798), .B(n5789), .Y(n5788) );
  BUFX3 U17088 ( .A(n11497), .Y(M3_mult_x_15_b_17_) );
  INVXL U17089 ( .A(n18080), .Y(n4733) );
  INVXL U17090 ( .A(n4733), .Y(n4734) );
  INVXL U17091 ( .A(n6408), .Y(n4735) );
  INVXL U17092 ( .A(n4735), .Y(n4736) );
  INVXL U17093 ( .A(n6611), .Y(n4737) );
  INVX1 U17094 ( .A(n4737), .Y(n4738) );
  OAI22X1 U17095 ( .A0(n9963), .A1(n9595), .B0(n9441), .B1(n3180), .Y(n9594)
         );
  BUFX4 U17096 ( .A(n9694), .Y(n9963) );
  OAI22X1 U17097 ( .A0(n9963), .A1(n9844), .B0(n9962), .B1(n3180), .Y(n9958)
         );
  INVXL U17098 ( .A(n12337), .Y(n4741) );
  INVXL U17099 ( .A(n4741), .Y(n4742) );
  OAI22X1 U17100 ( .A0(n14208), .A1(n14197), .B0(n13281), .B1(n14198), .Y(
        n13327) );
  OAI22X1 U17101 ( .A0(n6191), .A1(n14290), .B0(n13511), .B1(n14298), .Y(
        n13551) );
  OAI22X1 U17102 ( .A0(n16638), .A1(n16462), .B0(n16396), .B1(n16475), .Y(
        n16461) );
  XNOR2X1 U17103 ( .A(M5_mult_x_15_n1), .B(n3198), .Y(n16396) );
  XNOR2X1 U17104 ( .A(M4_a_1_), .B(M3_mult_x_15_b_21_), .Y(n17604) );
  NOR2X1 U17105 ( .A(n4581), .B(n6271), .Y(n24024) );
  XOR2XL U17106 ( .A(n22881), .B(n3053), .Y(M6_mult_x_15_n1177) );
  OAI222X1 U17107 ( .A0(n26540), .A1(n23884), .B0(n3121), .B1(n24129), .C0(
        n4586), .C1(n24515), .Y(n2609) );
  AOI22X2 U17108 ( .A0(n23741), .A1(n19104), .B0(n3128), .B1(n23521), .Y(
        n25483) );
  CMPR22X1 U17109 ( .A(n23776), .B(n23775), .CO(n20799), .S(n23777) );
  CMPR22X1 U17110 ( .A(n20791), .B(n20790), .CO(n23775), .S(n20792) );
  ADDHXL U17111 ( .A(n16642), .B(n16641), .CO(n16643), .S(n16634) );
  OAI22X1 U17112 ( .A0(n10295), .A1(n10325), .B0(n10326), .B1(n9799), .Y(n9818) );
  NAND2X2 U17113 ( .A(n9205), .B(n10326), .Y(n10325) );
  INVXL U17114 ( .A(n9957), .Y(n4743) );
  INVXL U17115 ( .A(n4743), .Y(n4744) );
  INVXL U17116 ( .A(n11817), .Y(n4745) );
  OAI22X1 U17117 ( .A0(n12598), .A1(n12225), .B0(n12342), .B1(n12224), .Y(
        n12336) );
  OAI22X1 U17118 ( .A0(n13328), .A1(n3181), .B0(n13282), .B1(n13532), .Y(
        n13326) );
  ADDHXL U17119 ( .A(n13499), .B(n13498), .CO(n13528), .S(n13475) );
  XNOR2XL U17120 ( .A(M0_b_9_), .B(n21054), .Y(n6501) );
  OAI22X1 U17121 ( .A0(n6524), .A1(n7094), .B0(n7093), .B1(n6523), .Y(n6690)
         );
  INVXL U17122 ( .A(n9238), .Y(n4747) );
  INVXL U17123 ( .A(n4747), .Y(n4748) );
  ADDFX2 U17124 ( .A(n9358), .B(n9357), .CI(n9356), .CO(n9457), .S(n9352) );
  ADDFX2 U17125 ( .A(n9749), .B(n9748), .CI(n9747), .CO(n9761), .S(n9788) );
  ADDFX2 U17126 ( .A(n11661), .B(n11660), .CI(n11659), .CO(n11693), .S(n11735)
         );
  ADDFX2 U17127 ( .A(n11777), .B(n11776), .CI(n11775), .CO(n11874), .S(n11771)
         );
  OAI22X1 U17128 ( .A0(n12352), .A1(n12034), .B0(n12222), .B1(n12033), .Y(
        n12057) );
  ADDFX2 U17129 ( .A(n16386), .B(n16385), .CI(n16384), .CO(n16395), .S(n16457)
         );
  OAI22X1 U17130 ( .A0(n18107), .A1(n17517), .B0(n17902), .B1(n17505), .Y(
        n17532) );
  INVXL U17131 ( .A(n17585), .Y(n4749) );
  INVX1 U17132 ( .A(n4749), .Y(n4750) );
  XOR2X1 U17133 ( .A(n11834), .B(n4926), .Y(n4925) );
  XNOR2X1 U17134 ( .A(n7286), .B(M0_b_13_), .Y(n6781) );
  OAI21X1 U17135 ( .A0(n6274), .A1(n26222), .B0(n6265), .Y(M0_b_13_) );
  NOR2X1 U17136 ( .A(n24856), .B(n23200), .Y(n24492) );
  CLKINVX3 U17137 ( .A(n14683), .Y(n4752) );
  OAI222X1 U17138 ( .A0(n6184), .A1(n11483), .B0(n25901), .B1(n25813), .C0(
        n15940), .C1(n23991), .Y(n11493) );
  XOR2X1 U17139 ( .A(n17776), .B(n4885), .Y(n4884) );
  OAI22X1 U17140 ( .A0(n18111), .A1(n17743), .B0(n18504), .B1(n17791), .Y(
        n17776) );
  INVX4 U17141 ( .A(n3118), .Y(n25292) );
  BUFX3 U17142 ( .A(n12523), .Y(n12595) );
  INVXL U17143 ( .A(n6793), .Y(n4755) );
  INVX1 U17144 ( .A(n4755), .Y(n4756) );
  OAI22X1 U17145 ( .A0(n10300), .A1(n10541), .B0(n10330), .B1(n3174), .Y(
        n10347) );
  OAI22X1 U17146 ( .A0(n10300), .A1(n3174), .B0(n10541), .B1(n10161), .Y(
        n10306) );
  INVXL U17147 ( .A(n6535), .Y(n4757) );
  INVXL U17148 ( .A(n4757), .Y(n4758) );
  INVXL U17149 ( .A(n6650), .Y(n4759) );
  INVXL U17150 ( .A(n4759), .Y(n4760) );
  OAI22X1 U17151 ( .A0(n6554), .A1(n7093), .B0(n6616), .B1(n7094), .Y(n6627)
         );
  OAI22X1 U17152 ( .A0(n6554), .A1(n7094), .B0(n7093), .B1(n6553), .Y(n6558)
         );
  OAI22X1 U17153 ( .A0(n7093), .A1(n6833), .B0(n6919), .B1(n7094), .Y(n6917)
         );
  ADDFX2 U17154 ( .A(n9213), .B(n9212), .CI(n9211), .CO(n9333), .S(n9289) );
  OAI22X1 U17155 ( .A0(n10541), .A1(n9266), .B0(n3174), .B1(n9210), .Y(n9212)
         );
  ADDFX2 U17156 ( .A(n10165), .B(n10164), .CI(n10163), .CO(n10294), .S(n10150)
         );
  OAI22X1 U17157 ( .A0(n10541), .A1(n9580), .B0(n10329), .B1(n10161), .Y(
        n10164) );
  OAI22X1 U17158 ( .A0(n10660), .A1(n10514), .B0(n3178), .B1(n10539), .Y(
        n10492) );
  OAI22X1 U17159 ( .A0(n12635), .A1(n12013), .B0(n12513), .B1(n11993), .Y(
        n12053) );
  XNOR2XL U17160 ( .A(n12519), .B(n3197), .Y(n11993) );
  OAI22XL U17161 ( .A0(n12598), .A1(n12219), .B0(n12342), .B1(n12343), .Y(
        n12345) );
  OAI22X1 U17162 ( .A0(n12293), .A1(n12255), .B0(n12245), .B1(n12338), .Y(
        n12258) );
  BUFX3 U17163 ( .A(n4775), .Y(n12338) );
  OAI22XL U17164 ( .A0(n13482), .A1(n13790), .B0(n13538), .B1(n13721), .Y(
        n13526) );
  ADDFX2 U17165 ( .A(n13554), .B(n13553), .CI(n13552), .CO(n13634), .S(n13569)
         );
  OAI22XL U17166 ( .A0(n13564), .A1(n3181), .B0(n13533), .B1(n13532), .Y(
        n13553) );
  INVXL U17167 ( .A(n13671), .Y(n4761) );
  INVXL U17168 ( .A(n4761), .Y(n4762) );
  OAI22X1 U17169 ( .A0(n13836), .A1(n14291), .B0(n13780), .B1(n6191), .Y(
        n13858) );
  OAI22X1 U17170 ( .A0(n14024), .A1(n6191), .B0(n14047), .B1(n14298), .Y(
        n14049) );
  OAI22X1 U17171 ( .A0(n2993), .A1(n14195), .B0(n14289), .B1(n14236), .Y(
        n14151) );
  ADDFX2 U17172 ( .A(n16316), .B(n16315), .CI(n16314), .CO(n16991), .S(n16301)
         );
  INVXL U17173 ( .A(n16365), .Y(n4763) );
  INVXL U17174 ( .A(n4763), .Y(n4764) );
  OAI22X1 U17175 ( .A0(n16638), .A1(n16576), .B0(n16575), .B1(n16475), .Y(
        n16579) );
  ADDFX2 U17176 ( .A(n17698), .B(n17697), .CI(n17696), .CO(n17684), .S(n18339)
         );
  OAI22XL U17177 ( .A0(n18177), .A1(n18139), .B0(n18129), .B1(n18223), .Y(
        n18144) );
  ADDFX2 U17178 ( .A(n5997), .B(n18647), .CI(n18646), .CO(n18656), .S(n18648)
         );
  CMPR22X1 U17179 ( .A(n20795), .B(n20794), .CO(n24274), .S(n20778) );
  INVXL U17180 ( .A(n23781), .Y(n4765) );
  INVXL U17181 ( .A(n4765), .Y(n4766) );
  NOR2X2 U17182 ( .A(n18675), .B(n18674), .Y(n18861) );
  OAI22X1 U17183 ( .A0(n21011), .A1(n21010), .B0(n3076), .B1(n21009), .Y(
        n24880) );
  XOR2XL U17184 ( .A(n17398), .B(n17397), .Y(n17192) );
  OAI22X1 U17185 ( .A0(n24858), .A1(n24857), .B0(n3074), .B1(n24856), .Y(
        n24951) );
  OAI21XL U17186 ( .A0(n23224), .A1(n23223), .B0(n3222), .Y(n23227) );
  CMPR22X1 U17187 ( .A(n9958), .B(n4744), .CO(n9995), .S(n9991) );
  CMPR22X1 U17188 ( .A(n4742), .B(n12336), .CO(n12369), .S(n12365) );
  OR2X2 U17189 ( .A(n24913), .B(n3121), .Y(n5599) );
  AOI2BB1X1 U17190 ( .A0N(n25783), .A1N(n3121), .B0(n4712), .Y(n25130) );
  AOI22X1 U17191 ( .A0(n20385), .A1(n23608), .B0(n25300), .B1(n23607), .Y(
        n23720) );
  INVX1 U17192 ( .A(n4770), .Y(n4771) );
  XOR2X1 U17193 ( .A(n17775), .B(n4884), .Y(n17793) );
  AOI22X1 U17194 ( .A0(n20385), .A1(n23616), .B0(n25300), .B1(n23615), .Y(
        n25323) );
  ADDFX2 U17195 ( .A(n7464), .B(n7463), .CI(n7462), .CO(n7505), .S(n7468) );
  OAI22X1 U17196 ( .A0(n10541), .A1(n9302), .B0(n3174), .B1(n9239), .Y(n9304)
         );
  INVXL U17197 ( .A(n11912), .Y(n4773) );
  INVX1 U17198 ( .A(n4773), .Y(n4774) );
  ADDFX2 U17199 ( .A(n12076), .B(n12075), .CI(n12074), .CO(n12091), .S(n12115)
         );
  OAI22XL U17200 ( .A0(n12618), .A1(n11743), .B0(n12119), .B1(n11723), .Y(
        n11797) );
  OAI22X1 U17201 ( .A0(n9551), .A1(n9207), .B0(n9838), .B1(n9220), .Y(n9279)
         );
  INVXL U17202 ( .A(n4775), .Y(n4776) );
  ADDFX2 U17203 ( .A(n9282), .B(n9281), .CI(n9280), .CO(n9336), .S(n9286) );
  XOR2X1 U17204 ( .A(n5995), .B(n12697), .Y(n12703) );
  CLKINVX3 U17205 ( .A(n13051), .Y(n13974) );
  ADDFX2 U17206 ( .A(n18022), .B(n18021), .CI(n18020), .CO(n18034), .S(n18055)
         );
  OAI22X1 U17207 ( .A0(n24724), .A1(n24723), .B0(n24722), .B1(n3074), .Y(
        n24808) );
  OAI211X4 U17208 ( .A0(n25903), .A1(n9087), .B0(n9061), .C0(n9060), .Y(
        M2_a_4_) );
  XOR2XL U17209 ( .A(n22612), .B(n3055), .Y(M6_mult_x_15_n1124) );
  XOR2XL U17210 ( .A(n22963), .B(n3055), .Y(M6_mult_x_15_n1123) );
  AOI22X1 U17211 ( .A0(n20385), .A1(n24785), .B0(n25300), .B1(n20852), .Y(
        n24741) );
  OAI21X1 U17212 ( .A0(n3073), .A1(n20431), .B0(n20430), .Y(n24785) );
  OAI22X1 U17213 ( .A0(n4592), .A1(n6314), .B0(n3046), .B1(n6313), .Y(n6338)
         );
  OAI22X1 U17214 ( .A0(n4592), .A1(n7564), .B0(n3046), .B1(n6398), .Y(n6435)
         );
  OAI222X4 U17215 ( .A0(n25895), .A1(n6274), .B0(n26287), .B1(n4583), .C0(
        n26025), .C1(n6266), .Y(M0_b_1_) );
  OAI222X4 U17216 ( .A0(n25896), .A1(n6274), .B0(n26027), .B1(n4583), .C0(
        n26256), .C1(n6266), .Y(M0_b_2_) );
  OAI21X2 U17217 ( .A0(n8482), .A1(n8167), .B0(n8166), .Y(n23858) );
  OAI21X2 U17218 ( .A0(n19564), .A1(n19301), .B0(n19300), .Y(n24341) );
  OAI21X2 U17219 ( .A0(n8482), .A1(n8171), .B0(n8170), .Y(n23810) );
  OAI21X2 U17220 ( .A0(n8482), .A1(n8169), .B0(n8168), .Y(n23816) );
  OAI21X2 U17221 ( .A0(n19566), .A1(n19299), .B0(n19298), .Y(n24072) );
  OAI222X4 U17222 ( .A0(n25991), .A1(n6274), .B0(n26260), .B1(n4583), .C0(
        n25888), .C1(n6266), .Y(M0_b_9_) );
  OAI21X1 U17223 ( .A0(n24315), .A1(n3024), .B0(n24313), .Y(n24314) );
  XOR2X1 U17224 ( .A(n5147), .B(n9677), .Y(n9719) );
  NOR2X2 U17225 ( .A(in_valid_t), .B(n3024), .Y(n25786) );
  CMPR22X1 U17226 ( .A(n14700), .B(n14713), .CO(n14461), .S(n24304) );
  OAI21X2 U17227 ( .A0(n19566), .A1(n19296), .B0(n19295), .Y(n24295) );
  OAI21X2 U17228 ( .A0(n19566), .A1(n19294), .B0(n19293), .Y(n24390) );
  NOR2X2 U17229 ( .A(n20379), .B(n9034), .Y(n23871) );
  AOI21X1 U17230 ( .A0(n9032), .A1(n9028), .B0(n9027), .Y(n9034) );
  XNOR2X2 U17231 ( .A(M5_a_12_), .B(n3203), .Y(n15996) );
  OAI222X4 U17232 ( .A0(n26518), .A1(n15942), .B0(n26279), .B1(n25813), .C0(
        n26034), .C1(n17167), .Y(M5_a_12_) );
  AOI21XL U17233 ( .A0(n24425), .A1(in_valid_d), .B0(n5561), .Y(n5560) );
  XOR2X1 U17234 ( .A(M3_mult_x_15_a_17_), .B(M3_a_16_), .Y(n5416) );
  AOI21XL U17235 ( .A0(n12696), .A1(n4918), .B0(M3_a_16_), .Y(
        M3_U3_U1_enc_tree_0__1__14_) );
  OAI22X1 U17236 ( .A0(n14249), .A1(n3019), .B0(n13362), .B1(n14250), .Y(
        n13366) );
  OAI22X1 U17237 ( .A0(n13403), .A1(n14249), .B0(n13422), .B1(n14250), .Y(
        n13435) );
  CLKINVX3 U17238 ( .A(n6208), .Y(n14250) );
  OAI21X1 U17239 ( .A0(n14833), .A1(n26189), .B0(n14843), .Y(n14951) );
  OAI222X1 U17240 ( .A0(n26539), .A1(n23884), .B0(n3121), .B1(n24132), .C0(
        n4584), .C1(n24536), .Y(n2607) );
  OAI22X1 U17241 ( .A0(n26141), .A1(n15942), .B0(n25915), .B1(n25813), .Y(
        n11482) );
  OAI21X1 U17242 ( .A0(n7148), .A1(n5124), .B0(n5115), .Y(n7181) );
  BUFX1 U17243 ( .A(n18147), .Y(n4799) );
  BUFX1 U17244 ( .A(n12262), .Y(n4800) );
  BUFX1 U17245 ( .A(n13090), .Y(n4801) );
  INVXL U17246 ( .A(n14937), .Y(n4802) );
  INVXL U17247 ( .A(n19340), .Y(n4803) );
  AOI22XL U17248 ( .A0(n25229), .A1(y12[18]), .B0(n14427), .B1(y10[18]), .Y(
        n9070) );
  NAND2X1 U17249 ( .A(n3132), .B(n20987), .Y(n5519) );
  NOR2X1 U17250 ( .A(n3146), .B(n3033), .Y(n23528) );
  NAND2X1 U17251 ( .A(n3132), .B(n23494), .Y(n5254) );
  OAI22X1 U17252 ( .A0(n12340), .A1(n12064), .B0(n12031), .B1(n12338), .Y(
        n12036) );
  NOR2X1 U17253 ( .A(n12985), .B(n12810), .Y(n12814) );
  CMPR22X1 U17254 ( .A(n25162), .B(n25159), .CO(n25131), .S(n25160) );
  CMPR22X1 U17255 ( .A(n25107), .B(n25106), .CO(n25159), .S(n25100) );
  CMPR22X1 U17256 ( .A(n25181), .B(n25178), .CO(n25106), .S(n25179) );
  CMPR22X1 U17257 ( .A(n23683), .B(n23682), .CO(n23849), .S(n7880) );
  CMPR22X1 U17258 ( .A(n23854), .B(n23853), .CO(n23682), .S(n23856) );
  CMPR22X1 U17259 ( .A(n24336), .B(n24335), .CO(n25183), .S(n24338) );
  CMPR22X1 U17260 ( .A(n24087), .B(n25804), .CO(n24335), .S(n24089) );
  CMPR22X1 U17261 ( .A(n24348), .B(n24347), .CO(n20794), .S(n24349) );
  CMPR22X1 U17262 ( .A(n20787), .B(n20786), .CO(n24347), .S(n20788) );
  OAI22X1 U17263 ( .A0(n10517), .A1(n5079), .B0(n10533), .B1(n9442), .Y(n9593)
         );
  BUFX1 U17264 ( .A(n16460), .Y(n4805) );
  OAI22X1 U17265 ( .A0(n6613), .A1(n6829), .B0(n6608), .B1(n6606), .Y(n6610)
         );
  ADDFX2 U17266 ( .A(n17712), .B(n17711), .CI(n17710), .CO(n18340), .S(n18366)
         );
  ADDFX2 U17267 ( .A(n16179), .B(n16178), .CI(n16177), .CO(n16198), .S(n16173)
         );
  OAI22X1 U17268 ( .A0(n16941), .A1(n16142), .B0(n16939), .B1(n16166), .Y(
        n16179) );
  OAI22XL U17269 ( .A0(n13727), .A1(n13971), .B0(n13777), .B1(n13972), .Y(
        n13796) );
  ADDFX2 U17270 ( .A(n6358), .B(n6357), .CI(n6356), .CO(n6769), .S(n6359) );
  ADDFX2 U17271 ( .A(n16492), .B(n16491), .CI(n16490), .CO(n16504), .S(n16556)
         );
  ADDFX2 U17272 ( .A(n12168), .B(n12167), .CI(n12166), .CO(n12159), .S(n12192)
         );
  NAND2X1 U17273 ( .A(n10615), .B(n10478), .Y(n5219) );
  XOR2X1 U17274 ( .A(n4931), .B(n21024), .Y(n24127) );
  XOR2X2 U17275 ( .A(n4993), .B(n20326), .Y(n24140) );
  OAI21XL U17276 ( .A0(n14533), .A1(n14487), .B0(n14486), .Y(n14496) );
  XOR2X1 U17277 ( .A(n5921), .B(n23478), .Y(n25590) );
  INVX1 U17278 ( .A(n14684), .Y(n20688) );
  AOI22X1 U17279 ( .A0(n4566), .A1(data[14]), .B0(n4579), .B1(w1[270]), .Y(
        n9080) );
  INVX1 U17280 ( .A(n20370), .Y(n5591) );
  XNOR2X1 U17281 ( .A(n10595), .B(n10594), .Y(n20711) );
  INVX1 U17282 ( .A(n19047), .Y(n5313) );
  NOR2X1 U17283 ( .A(n12489), .B(n12488), .Y(n12933) );
  INVX1 U17284 ( .A(n18972), .Y(n23733) );
  XOR2X1 U17285 ( .A(n20932), .B(n20931), .Y(n21049) );
  NOR2X1 U17286 ( .A(n20931), .B(n5750), .Y(n20920) );
  INVX1 U17287 ( .A(n18845), .Y(n5436) );
  OAI22X1 U17288 ( .A0(n12759), .A1(n12637), .B0(n12760), .B1(n12636), .Y(
        n12641) );
  OAI22X1 U17289 ( .A0(n10660), .A1(n10386), .B0(n3178), .B1(n10337), .Y(
        n10364) );
  OAI22X1 U17290 ( .A0(n10296), .A1(n9574), .B0(n10326), .B1(n10158), .Y(
        n10155) );
  OAI22X1 U17291 ( .A0(n16977), .A1(n16362), .B0(n3105), .B1(n16329), .Y(
        n16419) );
  OAI22X1 U17292 ( .A0(n7829), .A1(n7569), .B0(n7828), .B1(n25878), .Y(n7528)
         );
  OAI22XL U17293 ( .A0(n6613), .A1(n7088), .B0(n7146), .B1(n25867), .Y(n7157)
         );
  ADDFX2 U17294 ( .A(n6827), .B(n6826), .CI(n6825), .CO(n6950), .S(n6879) );
  OAI22X1 U17295 ( .A0(n7511), .A1(n6820), .B0(n7512), .B1(n6832), .Y(n6826)
         );
  OAI22X1 U17296 ( .A0(n9504), .A1(n9319), .B0(n10496), .B1(n9296), .Y(n9379)
         );
  OAI22X1 U17297 ( .A0(n10660), .A1(n9839), .B0(n3178), .B1(n10312), .Y(n9545)
         );
  OAI22X1 U17298 ( .A0(n10517), .A1(n9537), .B0(n10533), .B1(n9581), .Y(n9571)
         );
  ADDFX2 U17299 ( .A(n13562), .B(n13561), .CI(n13560), .CO(n13612), .S(n13557)
         );
  OAI22XL U17300 ( .A0(n13567), .A1(n14298), .B0(n13542), .B1(n6191), .Y(
        n13561) );
  ADDFX2 U17301 ( .A(n13958), .B(n13957), .CI(n13956), .CO(n14022), .S(n13978)
         );
  OAI22X1 U17302 ( .A0(n2993), .A1(n4567), .B0(n14356), .B1(n14118), .Y(n14061) );
  OAI22X1 U17303 ( .A0(n18522), .A1(n17969), .B0(n3195), .B1(n17968), .Y(
        n18003) );
  OAI22X1 U17304 ( .A0(n7829), .A1(n7164), .B0(n7828), .B1(n25882), .Y(n7100)
         );
  OAI22X1 U17305 ( .A0(n7535), .A1(n6311), .B0(n6751), .B1(n7460), .Y(n6754)
         );
  OAI22X1 U17306 ( .A0(n9694), .A1(n9441), .B0(n9405), .B1(n3180), .Y(n9597)
         );
  OAI22X1 U17307 ( .A0(n16941), .A1(n16409), .B0(n16939), .B1(n16346), .Y(
        n16413) );
  OAI22X1 U17308 ( .A0(n16941), .A1(n16513), .B0(n16939), .B1(n16468), .Y(
        n16500) );
  OAI22X1 U17309 ( .A0(n16941), .A1(n16539), .B0(n16939), .B1(n16538), .Y(
        n16706) );
  OAI22X1 U17310 ( .A0(n6489), .A1(n7511), .B0(n6542), .B1(n7512), .Y(n6544)
         );
  ADDFX2 U17311 ( .A(n6684), .B(n6683), .CI(n6682), .CO(n6699), .S(n6680) );
  ADDFX2 U17312 ( .A(n13377), .B(n13376), .CI(n13375), .CO(n13385), .S(n13382)
         );
  OAI22X1 U17313 ( .A0(n16638), .A1(n16603), .B0(n16593), .B1(n16475), .Y(
        n16607) );
  OAI22XL U17314 ( .A0(n12293), .A1(n12227), .B0(n12226), .B1(n12338), .Y(
        n12230) );
  OAI22X1 U17315 ( .A0(n13259), .A1(n14157), .B0(n13279), .B1(n14120), .Y(
        n13294) );
  OAI22X1 U17316 ( .A0(n9963), .A1(n9845), .B0(n9844), .B1(n3180), .Y(n9848)
         );
  ADDFX2 U17317 ( .A(n17615), .B(n17614), .CI(n17613), .CO(n17843), .S(n17642)
         );
  NOR2X1 U17318 ( .A(n20491), .B(n20473), .Y(n20502) );
  OAI22X1 U17319 ( .A0(n3031), .A1(n20392), .B0(n9005), .B1(n3071), .Y(n20491)
         );
  OAI21XL U17320 ( .A0(n17566), .A1(n5906), .B0(n17565), .Y(n5905) );
  XOR2XL U17321 ( .A(n22696), .B(n3053), .Y(M6_mult_x_15_n1173) );
  INVX1 U17322 ( .A(n20273), .Y(n20704) );
  INVX1 U17323 ( .A(n23706), .Y(n20663) );
  CMPR22X1 U17324 ( .A(n18088), .B(n18087), .CO(n18275), .S(n18217) );
  OAI22X1 U17325 ( .A0(n18083), .A1(n18428), .B0(n18429), .B1(n18068), .Y(
        n18087) );
  CMPR22X1 U17326 ( .A(n18221), .B(n18220), .CO(n18254), .S(n18250) );
  OAI22X1 U17327 ( .A0(n18111), .A1(n18110), .B0(n18504), .B1(n18109), .Y(
        n18220) );
  OAI22X1 U17328 ( .A0(n5466), .A1(n18177), .B0(n18223), .B1(n18225), .Y(
        n18221) );
  CMPR22X1 U17329 ( .A(n9658), .B(n9657), .CO(n9660), .S(n9678) );
  OAI22X1 U17330 ( .A0(n9504), .A1(n5202), .B0(n10496), .B1(n9632), .Y(n9657)
         );
  CMPR22X1 U17331 ( .A(n13366), .B(n13365), .CO(n13425), .S(n13378) );
  CMPR22X1 U17332 ( .A(n16683), .B(n16682), .CO(n16716), .S(n16712) );
  OAI22X1 U17333 ( .A0(n16942), .A1(n5729), .B0(n16943), .B1(n16574), .Y(
        n16682) );
  OAI22X1 U17334 ( .A0(n16638), .A1(n16575), .B0(n16685), .B1(n16475), .Y(
        n16683) );
  CMPR22X1 U17335 ( .A(n4740), .B(n12205), .CO(n12389), .S(n12333) );
  OAI22X1 U17336 ( .A0(n12597), .A1(n12522), .B0(n12595), .B1(n12187), .Y(
        n12205) );
  NAND2X1 U17337 ( .A(n17332), .B(n17331), .Y(n17333) );
  NAND2X1 U17338 ( .A(n10610), .B(n4611), .Y(n10611) );
  NAND2X1 U17339 ( .A(n17214), .B(n17213), .Y(n17215) );
  NAND2X1 U17340 ( .A(n18793), .B(n18831), .Y(n18794) );
  NAND2X1 U17341 ( .A(n3151), .B(n10206), .Y(n10207) );
  NAND2X1 U17342 ( .A(n7015), .B(n7014), .Y(n7016) );
  XOR2X1 U17343 ( .A(n5712), .B(n17234), .Y(n20744) );
  XOR2X2 U17344 ( .A(n5660), .B(n4679), .Y(n20926) );
  NAND2X1 U17345 ( .A(n17211), .B(n17229), .Y(n17212) );
  XOR2X2 U17346 ( .A(n13210), .B(n5163), .Y(n13235) );
  NOR2X2 U17347 ( .A(n10279), .B(n10283), .Y(n10197) );
  NOR2X1 U17348 ( .A(n10118), .B(n10117), .Y(n10279) );
  CMPR22X1 U17349 ( .A(n24110), .B(n24109), .CO(n25123), .S(n24111) );
  CMPR22X1 U17350 ( .A(n24275), .B(n24274), .CO(n24109), .S(n24276) );
  OAI22X1 U17351 ( .A0(n13555), .A1(n14282), .B0(n13621), .B1(n14251), .Y(
        n13598) );
  OAI22X1 U17352 ( .A0(n13737), .A1(n14282), .B0(n13778), .B1(n14251), .Y(
        n13798) );
  ADDFX2 U17353 ( .A(n16068), .B(n16067), .CI(n16066), .CO(n16096), .S(n16792)
         );
  ADDFX2 U17354 ( .A(n13574), .B(n13573), .CI(n13572), .CO(n13641), .S(n13558)
         );
  OAI22X2 U17355 ( .A0(n17937), .A1(n17973), .B0(n18168), .B1(n17936), .Y(
        n17977) );
  ADDFX2 U17356 ( .A(n16710), .B(n16709), .CI(n16708), .CO(n16740), .S(n16719)
         );
  ADDFX2 U17357 ( .A(n6405), .B(n6404), .CI(n6403), .CO(n6401), .S(n6448) );
  BUFX3 U17358 ( .A(M1_a_5_), .Y(n13919) );
  CLKINVX3 U17359 ( .A(n6299), .Y(n7615) );
  OAI21X2 U17360 ( .A0(n7382), .A1(n26010), .B0(n6280), .Y(n6299) );
  NOR2X2 U17361 ( .A(n14503), .B(n14346), .Y(n14673) );
  CMPR22X1 U17362 ( .A(n25099), .B(n25098), .CO(n25178), .S(n24361) );
  CMPR22X1 U17363 ( .A(n24360), .B(n24359), .CO(n25098), .S(n23646) );
  CMPR22X1 U17364 ( .A(n23822), .B(n23821), .CO(n23853), .S(n23824) );
  CMPR22X1 U17365 ( .A(n23782), .B(n4766), .CO(n23821), .S(n23783) );
  OAI22XL U17366 ( .A0(n12635), .A1(n12102), .B0(n12513), .B1(n12066), .Y(
        n12107) );
  INVX1 U17367 ( .A(n10713), .Y(n5479) );
  NAND2BX1 U17368 ( .AN(n17740), .B(n5885), .Y(n5884) );
  OAI2BB1X1 U17369 ( .A0N(n17740), .A1N(n5887), .B0(n5883), .Y(n17794) );
  OAI22X1 U17370 ( .A0(n18522), .A1(n17734), .B0(n3195), .B1(n17741), .Y(
        n17740) );
  NAND2X1 U17371 ( .A(n7672), .B(n7779), .Y(n7815) );
  XOR2X1 U17372 ( .A(n17729), .B(n5796), .Y(n17768) );
  XOR3X2 U17373 ( .A(n13605), .B(n6053), .C(n13732), .Y(n5215) );
  XNOR2X1 U17374 ( .A(n9797), .B(n5188), .Y(n5187) );
  OAI22X1 U17375 ( .A0(n9983), .A1(n9785), .B0(n9981), .B1(n9754), .Y(n5188)
         );
  AOI21X1 U17376 ( .A0(n10642), .A1(n10641), .B0(n10640), .Y(n5249) );
  OAI2BB1X1 U17377 ( .A0N(n5300), .A1N(n9477), .B0(n5299), .Y(n9497) );
  XOR2XL U17378 ( .A(M4_a_18_), .B(M4_a_19_), .Y(n17494) );
  ADDFX2 U17379 ( .A(n12558), .B(n12557), .CI(n12556), .CO(n12582), .S(n12551)
         );
  ADDFX2 U17380 ( .A(n9500), .B(n9499), .CI(n9498), .CO(n9554), .S(n9496) );
  ADDFX2 U17381 ( .A(n9777), .B(n9776), .CI(n9775), .CO(n9768), .S(n9804) );
  NAND2X1 U17382 ( .A(n12782), .B(n12781), .Y(n12867) );
  OAI22XL U17383 ( .A0(n9979), .A1(n9786), .B0(n9977), .B1(n9755), .Y(n9796)
         );
  XOR2X1 U17384 ( .A(n16971), .B(n5671), .Y(n16992) );
  XOR2X1 U17385 ( .A(n5530), .B(n9423), .Y(n10069) );
  XNOR3X2 U17386 ( .A(n4914), .B(n12644), .C(n12643), .Y(n12658) );
  OAI2BB1X1 U17387 ( .A0N(n12698), .A1N(n5996), .B0(n5993), .Y(n12720) );
  OAI22X1 U17388 ( .A0(n15817), .A1(n15816), .B0(n15815), .B1(n3076), .Y(
        n24771) );
  AOI21X2 U17389 ( .A0(n14522), .A1(n14526), .B0(n14321), .Y(n5392) );
  NOR2X1 U17390 ( .A(n20617), .B(n20616), .Y(n5574) );
  INVX1 U17391 ( .A(n24044), .Y(n6107) );
  OAI211X4 U17392 ( .A0(n25900), .A1(n9087), .B0(n9052), .C0(n9051), .Y(
        M2_a_2_) );
  XOR2X2 U17393 ( .A(n23176), .B(n23177), .Y(n8823) );
  AOI21XL U17394 ( .A0(n24993), .A1(n20182), .B0(n24992), .Y(n24996) );
  NOR2X1 U17395 ( .A(n20181), .B(n20182), .Y(n20246) );
  OAI22X1 U17396 ( .A0(n13481), .A1(n14029), .B0(n13421), .B1(n14044), .Y(
        n13480) );
  OAI22X1 U17397 ( .A0(n13155), .A1(n14029), .B0(n13043), .B1(n14044), .Y(
        n13163) );
  NOR2X1 U17398 ( .A(n15940), .B(n23994), .Y(n5433) );
  OAI22X1 U17399 ( .A0(n12995), .A1(n12271), .B0(n12535), .B1(
        M3_mult_x_15_b_1_), .Y(n11646) );
  OAI22X1 U17400 ( .A0(n12535), .A1(n3108), .B0(n12995), .B1(n3049), .Y(n11881) );
  OAI22X1 U17401 ( .A0(n12535), .A1(n3197), .B0(n12995), .B1(
        M3_mult_x_15_n1682), .Y(n11953) );
  OAI22X1 U17402 ( .A0(n12535), .A1(M3_mult_x_15_b_9_), .B0(n12995), .B1(
        n16884), .Y(n12621) );
  OAI22X1 U17403 ( .A0(n3190), .A1(n12535), .B0(n12561), .B1(n12521), .Y(
        n12591) );
  NAND3X2 U17404 ( .A(n11551), .B(n11550), .C(n11549), .Y(n18767) );
  XOR2XL U17405 ( .A(n22864), .B(n3054), .Y(M6_mult_x_15_n1146) );
  XOR2XL U17406 ( .A(n22957), .B(n3054), .Y(M6_mult_x_15_n1148) );
  XOR2XL U17407 ( .A(n22837), .B(n3055), .Y(M6_mult_x_15_n1119) );
  XOR2XL U17408 ( .A(n22803), .B(n3055), .Y(M6_mult_x_15_n1118) );
  XOR2XL U17409 ( .A(n22654), .B(n3056), .Y(M6_mult_x_15_n1091) );
  XOR2XL U17410 ( .A(n22862), .B(n3056), .Y(M6_mult_x_15_n1094) );
  INVX1 U17411 ( .A(n12020), .Y(n5780) );
  XNOR2X1 U17412 ( .A(n3022), .B(n3198), .Y(n16871) );
  NOR2X1 U17413 ( .A(n17371), .B(n17374), .Y(n17377) );
  NOR2BX1 U17414 ( .AN(n6944), .B(n7512), .Y(n6499) );
  NOR2X1 U17415 ( .A(n17387), .B(n17391), .Y(n17360) );
  INVX1 U17416 ( .A(n19048), .Y(n5208) );
  XOR2XL U17417 ( .A(n22572), .B(n3119), .Y(M6_mult_x_15_n1037) );
  XOR2XL U17418 ( .A(n22598), .B(n3119), .Y(M6_mult_x_15_n1038) );
  XOR2XL U17419 ( .A(n22634), .B(n3119), .Y(n22635) );
  INVX1 U17420 ( .A(n19912), .Y(n19992) );
  OAI22X1 U17421 ( .A0(n4569), .A1(n10388), .B0(n10403), .B1(n9695), .Y(n9722)
         );
  OAI21XL U17422 ( .A0(n25851), .A1(n3024), .B0(n25817), .Y(n25818) );
  OAI21XL U17423 ( .A0(n24449), .A1(n3024), .B0(n24394), .Y(n24395) );
  NOR2X2 U17424 ( .A(n9033), .B(n9034), .Y(n23873) );
  NOR2X2 U17425 ( .A(n24069), .B(n24071), .Y(n24436) );
  NOR2X2 U17426 ( .A(n23958), .B(n23959), .Y(n24430) );
  AOI21XL U17427 ( .A0(n19954), .A1(n19952), .B0(n3164), .Y(n19953) );
  AOI21XL U17428 ( .A0(n19926), .A1(n19952), .B0(n3164), .Y(n19925) );
  AOI21XL U17429 ( .A0(n19931), .A1(n19952), .B0(n3164), .Y(n19930) );
  AOI21XL U17430 ( .A0(n19916), .A1(n19952), .B0(n3164), .Y(n19915) );
  OAI22X1 U17431 ( .A0(n13056), .A1(n13606), .B0(n13055), .B1(n3181), .Y(
        n13060) );
  NAND2X2 U17432 ( .A(n19654), .B(n19418), .Y(n19748) );
  NOR3X4 U17433 ( .A(n4768), .B(n23226), .C(n23225), .Y(n23415) );
  NAND3X1 U17434 ( .A(n24038), .B(n24039), .C(n25779), .Y(n25674) );
  NAND3X1 U17435 ( .A(n25780), .B(n25781), .C(n25779), .Y(n25819) );
  NAND3X1 U17436 ( .A(n24306), .B(n24307), .C(n25779), .Y(n25803) );
  NAND3X1 U17437 ( .A(n24282), .B(n24283), .C(n25779), .Y(n25170) );
  NAND3X1 U17438 ( .A(n24412), .B(n24413), .C(n25779), .Y(n25678) );
  NOR2X1 U17439 ( .A(n24626), .B(n25255), .Y(n24167) );
  OAI22X1 U17440 ( .A0(n16704), .A1(n3047), .B0(n5835), .B1(n16631), .Y(n16130) );
  OR2X2 U17441 ( .A(n16408), .B(n16704), .Y(n5860) );
  OAI22X1 U17442 ( .A0(n16704), .A1(n16380), .B0(n5835), .B1(n16116), .Y(
        n16430) );
  NAND2X2 U17443 ( .A(M4_a_1_), .B(n17962), .Y(n18226) );
  INVX1 U17444 ( .A(M4_a_0_), .Y(n17962) );
  CLKINVX3 U17445 ( .A(n23764), .Y(n24958) );
  OAI22XL U17446 ( .A0(n6991), .A1(n6481), .B0(n6602), .B1(n6490), .Y(n6498)
         );
  OAI2BB1X1 U17447 ( .A0N(n14081), .A1N(n14080), .B0(n25861), .Y(n14129) );
  OAI22X1 U17448 ( .A0(n4592), .A1(n7466), .B0(n3046), .B1(n7510), .Y(n7502)
         );
  OAI22X1 U17449 ( .A0(n4592), .A1(n7510), .B0(n3046), .B1(n7531), .Y(n7525)
         );
  AOI21XL U17450 ( .A0(n15536), .A1(n23955), .B0(n15573), .Y(n15535) );
  AOI21XL U17451 ( .A0(n15168), .A1(n23955), .B0(n15573), .Y(n15167) );
  AOI21XL U17452 ( .A0(n15221), .A1(n23955), .B0(n15573), .Y(n15220) );
  AOI222XL U17453 ( .A0(n23152), .A1(n11074), .B0(n23093), .B1(n3219), .C0(
        n23150), .C1(n11073), .Y(n22546) );
  AOI222XL U17454 ( .A0(n23152), .A1(n11062), .B0(n23093), .B1(n3217), .C0(
        n23150), .C1(n26493), .Y(n23134) );
  AOI222XL U17455 ( .A0(n23152), .A1(n3217), .B0(n23093), .B1(n23022), .C0(
        n23150), .C1(n11059), .Y(n22577) );
  AOI222XL U17456 ( .A0(n22928), .A1(n11073), .B0(n22700), .B1(n11063), .C0(
        n22927), .C1(n23109), .Y(n22627) );
  AOI222XL U17457 ( .A0(n22928), .A1(n11063), .B0(n22700), .B1(n23109), .C0(
        n22927), .C1(n11062), .Y(n22824) );
  AOI222XL U17458 ( .A0(n22928), .A1(n11062), .B0(n22700), .B1(n3217), .C0(
        n22927), .C1(n26493), .Y(n22853) );
  AOI222XL U17459 ( .A0(n22892), .A1(n3218), .B0(n22708), .B1(n23089), .C0(
        n22891), .C1(n11074), .Y(n22524) );
  AOI222XL U17460 ( .A0(n22892), .A1(n26493), .B0(n22708), .B1(n11059), .C0(
        n22891), .C1(n11058), .Y(n22831) );
  AOI222XL U17461 ( .A0(n22892), .A1(n3220), .B0(n22708), .B1(n22867), .C0(
        n22891), .C1(n10775), .Y(n22757) );
  AOI222XL U17462 ( .A0(n22892), .A1(n23151), .B0(n22708), .B1(n10789), .C0(
        n22891), .C1(n3220), .Y(n22874) );
  OAI21XL U17463 ( .A0(n9322), .A1(n9966), .B0(n6064), .Y(n9308) );
  OAI22X1 U17464 ( .A0(n9966), .A1(n9443), .B0(n10159), .B1(n9420), .Y(n9437)
         );
  OAI22X1 U17465 ( .A0(n12598), .A1(n11914), .B0(n12342), .B1(n11958), .Y(
        n11945) );
  OAI22X2 U17466 ( .A0(n13496), .A1(n14227), .B0(n13422), .B1(n14249), .Y(
        n13479) );
  CLKINVX3 U17467 ( .A(n6208), .Y(n14227) );
  OAI22X1 U17468 ( .A0(n10660), .A1(n10341), .B0(n10387), .B1(n3178), .Y(
        n10344) );
  XNOR2XL U17469 ( .A(n10494), .B(n10341), .Y(n9507) );
  XNOR2X1 U17470 ( .A(n10341), .B(M2_mult_x_15_a_1_), .Y(n5296) );
  BUFX3 U17471 ( .A(n7055), .Y(n4806) );
  OAI21XL U17472 ( .A0(n6274), .A1(n25894), .B0(n5579), .Y(n7055) );
  AOI2BB1X1 U17473 ( .A0N(n25687), .A1N(n4585), .B0(n4840), .Y(n20965) );
  AOI2BB1X1 U17474 ( .A0N(n23509), .A1N(n4583), .B0(n23508), .Y(n23510) );
  XOR2XL U17475 ( .A(n12716), .B(n6112), .Y(n12539) );
  XOR2XL U17476 ( .A(n12758), .B(n6112), .Y(n12713) );
  XOR2XL U17477 ( .A(n12265), .B(n6112), .Y(n11653) );
  XOR2X1 U17478 ( .A(n12594), .B(n6112), .Y(n11950) );
  XOR2X1 U17479 ( .A(n12732), .B(n6112), .Y(n12574) );
  XOR2X1 U17480 ( .A(n3204), .B(n6112), .Y(n11879) );
  XOR2X1 U17481 ( .A(n2980), .B(n6112), .Y(n11819) );
  XOR2X1 U17482 ( .A(n17073), .B(n16965), .Y(n16128) );
  XNOR2X1 U17483 ( .A(n17073), .B(M3_mult_x_15_b_21_), .Y(n17044) );
  XOR2XL U17484 ( .A(n3200), .B(n17073), .Y(n5096) );
  OAI22X1 U17485 ( .A0(n18541), .A1(n18042), .B0(n5893), .B1(n6129), .Y(n18061) );
  OAI22X1 U17486 ( .A0(n18541), .A1(n17882), .B0(n18539), .B1(n17862), .Y(
        n17916) );
  INVX1 U17487 ( .A(M4_mult_x_15_n1680), .Y(n18498) );
  XNOR2XL U17488 ( .A(n12233), .B(M4_mult_x_15_n1680), .Y(n12073) );
  OAI22X1 U17489 ( .A0(n18721), .A1(M3_mult_x_15_b_9_), .B0(n17512), .B1(
        M4_mult_x_15_n1680), .Y(n18525) );
  XNOR2XL U17490 ( .A(n18150), .B(M4_mult_x_15_n1680), .Y(n18005) );
  XNOR2X1 U17491 ( .A(n25884), .B(M4_mult_x_15_n1680), .Y(n11651) );
  XNOR2XL U17492 ( .A(n25883), .B(M4_mult_x_15_n1680), .Y(n17777) );
  XNOR2XL U17493 ( .A(n18503), .B(M4_mult_x_15_n1680), .Y(n17893) );
  XNOR2XL U17494 ( .A(n18118), .B(M4_mult_x_15_n1680), .Y(n17943) );
  XNOR2XL U17495 ( .A(n18006), .B(M4_mult_x_15_n1680), .Y(n18224) );
  XNOR2XL U17496 ( .A(n18500), .B(M4_mult_x_15_n1680), .Y(n17707) );
  XNOR2X1 U17497 ( .A(n18468), .B(M4_mult_x_15_n1680), .Y(n17518) );
  XNOR2XL U17498 ( .A(n18604), .B(M4_mult_x_15_n1680), .Y(n17506) );
  INVX8 U17499 ( .A(n25059), .Y(n25822) );
  CLKINVX3 U17500 ( .A(n5202), .Y(n4808) );
  NAND2X1 U17501 ( .A(n23707), .B(n5389), .Y(n20687) );
  OAI22XL U17502 ( .A0(n13932), .A1(n3173), .B0(n13874), .B1(n14080), .Y(
        n13931) );
  INVX1 U17503 ( .A(n14686), .Y(n23648) );
  AOI22X2 U17504 ( .A0(n20690), .A1(n3081), .B0(n4267), .B1(n23882), .Y(n24936) );
  XOR2X2 U17505 ( .A(n3212), .B(n4794), .Y(n5676) );
  INVX1 U17506 ( .A(n5100), .Y(n4809) );
  INVX1 U17507 ( .A(n14533), .Y(n14674) );
  CMPR22X1 U17508 ( .A(n11818), .B(n4746), .CO(n11841), .S(n12449) );
  NOR2X1 U17509 ( .A(n25767), .B(n25900), .Y(n6156) );
  OR2X2 U17510 ( .A(n16889), .B(n17092), .Y(n5827) );
  XNOR2X1 U17511 ( .A(M2_mult_x_15_n43), .B(n10335), .Y(n9549) );
  AOI22XL U17512 ( .A0(n25229), .A1(y12[20]), .B0(n14427), .B1(y10[20]), .Y(
        n9082) );
  CLKINVX3 U17513 ( .A(n23807), .Y(n5587) );
  OAI21X1 U17514 ( .A0(n18328), .A1(n18327), .B0(n18326), .Y(n18329) );
  XNOR2X1 U17515 ( .A(n25861), .B(n25865), .Y(n13283) );
  NAND2X1 U17516 ( .A(n5537), .B(n5535), .Y(n5534) );
  XNOR2X1 U17517 ( .A(n9904), .B(n10538), .Y(n9384) );
  OAI22X1 U17518 ( .A0(n6923), .A1(n7695), .B0(n6842), .B1(n5124), .Y(n6946)
         );
  NAND2X1 U17519 ( .A(n3132), .B(n20272), .Y(n20274) );
  NAND2BXL U17520 ( .AN(n9960), .B(n4808), .Y(n9632) );
  ADDFHX2 U17521 ( .A(n13756), .B(n13755), .CI(n13754), .CO(n13801), .S(n13818) );
  OAI21XL U17522 ( .A0(n19707), .A1(n20034), .B0(n19706), .Y(n20018) );
  INVX1 U17523 ( .A(M2_a_0_), .Y(n9781) );
  NAND2X1 U17524 ( .A(n14728), .B(n23744), .Y(n14729) );
  XNOR2X1 U17525 ( .A(n20025), .B(n20024), .Y(n20177) );
  CLKINVX3 U17526 ( .A(n19730), .Y(n19747) );
  NOR2X1 U17527 ( .A(n24391), .B(n20121), .Y(n20119) );
  XNOR2X1 U17528 ( .A(n14118), .B(n25862), .Y(n13700) );
  XNOR2X1 U17529 ( .A(n14357), .B(n13605), .Y(n13607) );
  AOI21X1 U17530 ( .A0(n6066), .A1(n14633), .B0(n14615), .Y(n14616) );
  XOR2X2 U17531 ( .A(n10222), .B(n4613), .Y(n19074) );
  INVX1 U17532 ( .A(n20099), .Y(n20101) );
  INVX1 U17533 ( .A(n20265), .Y(n25485) );
  AOI21X1 U17534 ( .A0(n19402), .A1(n19401), .B0(n19400), .Y(n19423) );
  NAND3BX2 U17535 ( .AN(n5182), .B(n9076), .C(n9075), .Y(M2_a_16_) );
  OAI21XL U17536 ( .A0(n25483), .A1(n3059), .B0(n20266), .Y(n20267) );
  AOI2BB1X1 U17537 ( .A0N(n3168), .A1N(n7445), .B0(n7444), .Y(n5126) );
  NOR2X2 U17538 ( .A(n5655), .B(n16506), .Y(n5654) );
  OAI22X1 U17539 ( .A0(n7287), .A1(n6831), .B0(n6929), .B1(n7288), .Y(n6927)
         );
  OAI21XL U17540 ( .A0(n8625), .A1(n8905), .B0(n8624), .Y(n8889) );
  XNOR2X1 U17541 ( .A(M2_mult_x_15_n43), .B(n9901), .Y(n9651) );
  XNOR2X1 U17542 ( .A(M2_mult_x_15_n43), .B(M2_mult_x_15_n1669), .Y(n10333) );
  OAI21XL U17543 ( .A0(n9287), .A1(n9288), .B0(n9286), .Y(n4816) );
  XOR3X2 U17544 ( .A(n9288), .B(n9286), .C(n9287), .Y(n9293) );
  NAND3BX2 U17545 ( .AN(n19100), .B(n3132), .C(n5191), .Y(n5190) );
  AOI22X1 U17546 ( .A0(n5336), .A1(n20938), .B0(n20933), .B1(n3136), .Y(n24248) );
  INVXL U17547 ( .A(n17332), .Y(n17114) );
  OAI22X1 U17548 ( .A0(n16977), .A1(n16976), .B0(n3105), .B1(n16975), .Y(
        n16984) );
  OAI21X1 U17549 ( .A0(n10185), .A1(n10243), .B0(n10184), .Y(n10189) );
  XNOR2X1 U17550 ( .A(n9904), .B(M2_mult_x_15_n1669), .Y(n9253) );
  NAND2X1 U17551 ( .A(n18406), .B(n18405), .Y(n18909) );
  AOI21XL U17552 ( .A0(n25754), .A1(n25170), .B0(n25169), .Y(n2351) );
  OAI21X1 U17553 ( .A0(n18880), .A1(n18925), .B0(n18879), .Y(n18885) );
  XNOR2X1 U17554 ( .A(n17039), .B(n3197), .Y(n15966) );
  OAI22X1 U17555 ( .A0(n17092), .A1(n16004), .B0(n16317), .B1(n16003), .Y(
        n16027) );
  AOI2BB1X1 U17556 ( .A0N(n24783), .A1N(n4586), .B0(n4823), .Y(n20775) );
  NAND3X4 U17557 ( .A(n4825), .B(n6149), .C(n6148), .Y(M4_mult_x_15_n1680) );
  INVX1 U17558 ( .A(n23770), .Y(n24475) );
  NAND2X1 U17559 ( .A(n6715), .B(n6714), .Y(n6716) );
  XNOR2X1 U17560 ( .A(n18872), .B(n18871), .Y(n23513) );
  INVX4 U17561 ( .A(n18918), .Y(n18925) );
  BUFX8 U17562 ( .A(n9164), .Y(n4826) );
  ADDFHX2 U17563 ( .A(n13439), .B(n13438), .CI(n13437), .CO(n13504), .S(n13455) );
  ADDFX2 U17564 ( .A(n13398), .B(n13397), .CI(n13396), .CO(n13442), .S(n13406)
         );
  NOR2X2 U17565 ( .A(n5468), .B(n4659), .Y(n5481) );
  OAI21X1 U17566 ( .A0(n7438), .A1(n7448), .B0(n7439), .Y(n7270) );
  NOR2X1 U17567 ( .A(n23709), .B(n23708), .Y(n23710) );
  NOR2X2 U17568 ( .A(n7360), .B(n7365), .Y(n7019) );
  NAND2X1 U17569 ( .A(n20700), .B(n23734), .Y(n5799) );
  OAI22X1 U17570 ( .A0(n18541), .A1(n17901), .B0(n5893), .B1(n17882), .Y(
        n17886) );
  INVX1 U17571 ( .A(n18866), .Y(n18896) );
  XOR2X1 U17572 ( .A(n11785), .B(n11784), .Y(n4865) );
  AOI21X1 U17573 ( .A0(n6733), .A1(y10[4]), .B0(n25142), .Y(n6261) );
  OAI21X2 U17574 ( .A0(n7382), .A1(n26001), .B0(n6261), .Y(M0_a_4_) );
  NAND2X1 U17575 ( .A(n23744), .B(n19091), .Y(n19093) );
  XNOR2X1 U17576 ( .A(n25864), .B(n25863), .Y(n14158) );
  XNOR2X1 U17577 ( .A(n12233), .B(n3201), .Y(n11721) );
  NAND2BX1 U17578 ( .AN(n13348), .B(n5024), .Y(n13350) );
  OAI21XL U17579 ( .A0(n17305), .A1(n17219), .B0(n17218), .Y(n17224) );
  XOR2X2 U17580 ( .A(n10189), .B(n4614), .Y(n17484) );
  NAND2X1 U17581 ( .A(n16849), .B(n16848), .Y(n17208) );
  AOI21X2 U17582 ( .A0(n11536), .A1(n4723), .B0(n5239), .Y(n5203) );
  NAND2X1 U17583 ( .A(n5701), .B(n5707), .Y(mul5_out[12]) );
  OAI22X1 U17584 ( .A0(n17092), .A1(n15972), .B0(n16317), .B1(n16004), .Y(
        n15985) );
  NAND2X1 U17585 ( .A(n17450), .B(n17452), .Y(n17420) );
  OAI22X1 U17586 ( .A0(n17092), .A1(n16184), .B0(n16317), .B1(n16203), .Y(
        n16217) );
  AOI22X1 U17587 ( .A0(n25229), .A1(y12[8]), .B0(n14427), .B1(y10[8]), .Y(
        n9092) );
  XOR3X2 U17588 ( .A(n14108), .B(n14111), .C(n14110), .Y(n14113) );
  AOI21X4 U17589 ( .A0(n6066), .A1(n5210), .B0(n13991), .Y(n14623) );
  NAND2X1 U17590 ( .A(n3132), .B(n20811), .Y(n20813) );
  OR2X2 U17591 ( .A(n18320), .B(n18319), .Y(n17985) );
  XOR2X2 U17592 ( .A(n7787), .B(n4641), .Y(n20759) );
  XNOR2X2 U17593 ( .A(n7720), .B(n7719), .Y(n20618) );
  OAI22X1 U17594 ( .A0(n6845), .A1(n6470), .B0(n6450), .B1(n6843), .Y(n6538)
         );
  BUFX3 U17595 ( .A(n17902), .Y(n18235) );
  OAI22XL U17596 ( .A0(n9983), .A1(n9730), .B0(n9906), .B1(n9706), .Y(n9746)
         );
  ADDFHX4 U17597 ( .A(n16437), .B(n16436), .CI(n16435), .CO(n16832), .S(n16433) );
  AOI21X2 U17598 ( .A0(n4875), .A1(data[49]), .B0(n5418), .Y(n5417) );
  XNOR2X1 U17599 ( .A(n18118), .B(M3_mult_x_15_b_21_), .Y(n17620) );
  OAI22X1 U17600 ( .A0(n6991), .A1(n6367), .B0(n6990), .B1(n6302), .Y(n6369)
         );
  OAI22X1 U17601 ( .A0(n4642), .A1(n7025), .B0(n7047), .B1(n7712), .Y(n7063)
         );
  ADDFHX2 U17602 ( .A(n16826), .B(n16825), .CI(n16824), .CO(n16846), .S(n16845) );
  NAND2XL U17603 ( .A(n9684), .B(n9686), .Y(n4830) );
  XOR3X2 U17604 ( .A(n9686), .B(n9684), .C(n9685), .Y(n9687) );
  CMPR22X1 U17605 ( .A(n6860), .B(n4804), .CO(n6939), .S(n6857) );
  ADDFHX1 U17606 ( .A(n16790), .B(n16789), .CI(n16788), .CO(n16805), .S(n16823) );
  NAND2X2 U17607 ( .A(n7004), .B(n7003), .Y(n7255) );
  OAI22X1 U17608 ( .A0(n17092), .A1(n16003), .B0(n16317), .B1(n15962), .Y(
        n15952) );
  CLKINVX8 U17609 ( .A(n7826), .Y(n7828) );
  NAND2X1 U17610 ( .A(n4834), .B(n4833), .Y(n17955) );
  XNOR3X2 U17611 ( .A(n17950), .B(n17951), .C(n4835), .Y(n17982) );
  INVX8 U17612 ( .A(n12751), .Y(n12758) );
  NAND2X1 U17613 ( .A(n21019), .B(n20315), .Y(n4983) );
  XOR2X2 U17614 ( .A(n4789), .B(M0_a_10_), .Y(n6275) );
  INVX1 U17615 ( .A(n17304), .Y(n17226) );
  XOR3X2 U17616 ( .A(n15995), .B(n15993), .C(n15994), .Y(n16083) );
  OAI22X1 U17617 ( .A0(n6991), .A1(n6775), .B0(n6990), .B1(n6835), .Y(n6867)
         );
  NAND3X1 U17618 ( .A(n5268), .B(n24189), .C(n5267), .Y(n5270) );
  OAI22X1 U17619 ( .A0(n18239), .A1(n17520), .B0(n18141), .B1(n17503), .Y(
        n17533) );
  OAI22X1 U17620 ( .A0(n17074), .A1(n16274), .B0(n16375), .B1(n16320), .Y(
        n16309) );
  INVX1 U17621 ( .A(n18948), .Y(n18939) );
  ADDFHX2 U17622 ( .A(n17847), .B(n17846), .CI(n17845), .CO(n17858), .S(n17855) );
  XOR2X1 U17623 ( .A(n4865), .B(n4863), .Y(n11788) );
  AOI21X1 U17624 ( .A0(n5990), .A1(n25796), .B0(n20843), .Y(n2285) );
  AOI22X1 U17625 ( .A0(n5480), .A1(sigma11[14]), .B0(in_valid_t), .B1(w2[46]), 
        .Y(n17473) );
  NOR2X1 U17626 ( .A(n6906), .B(n6905), .Y(n7360) );
  OAI22X1 U17627 ( .A0(n3102), .A1(n16219), .B0(n16332), .B1(n16289), .Y(
        n16236) );
  AOI21X1 U17628 ( .A0(n7364), .A1(n7012), .B0(n7011), .Y(n7017) );
  AOI21X1 U17629 ( .A0(n17462), .A1(n20353), .B0(n17461), .Y(n2284) );
  NAND2X1 U17630 ( .A(n3080), .B(n24206), .Y(n5514) );
  OAI22X1 U17631 ( .A0(n17092), .A1(n16978), .B0(n17099), .B1(n16875), .Y(
        n16945) );
  NAND2X2 U17632 ( .A(n14001), .B(n14594), .Y(n5278) );
  XOR2X2 U17633 ( .A(n17565), .B(n5908), .Y(n17573) );
  NOR2X1 U17634 ( .A(n18235), .B(n17504), .Y(n4847) );
  NOR2BX2 U17635 ( .AN(n12838), .B(n4891), .Y(n12846) );
  NOR2X4 U17636 ( .A(n7258), .B(n7259), .Y(n7308) );
  OAI22X1 U17637 ( .A0(n7511), .A1(n6964), .B0(n7512), .B1(n7051), .Y(n7033)
         );
  NOR2X2 U17638 ( .A(n5315), .B(n20810), .Y(n5314) );
  XNOR2XL U17639 ( .A(n3206), .B(M3_mult_x_15_b_13_), .Y(n17973) );
  XNOR2X4 U17640 ( .A(n5650), .B(n4682), .Y(n17464) );
  XNOR3X2 U17641 ( .A(n16077), .B(n6119), .C(n16076), .Y(n16078) );
  OAI22X1 U17642 ( .A0(n3102), .A1(n16088), .B0(n16332), .B1(n16009), .Y(
        n16068) );
  XOR2X2 U17643 ( .A(n4850), .B(n16416), .Y(n16453) );
  NOR2X2 U17644 ( .A(n5403), .B(n5402), .Y(n5966) );
  NAND2X1 U17645 ( .A(n17766), .B(n17765), .Y(n17806) );
  XNOR2X1 U17646 ( .A(n25883), .B(n3197), .Y(n17637) );
  NAND2X2 U17647 ( .A(n18675), .B(n18674), .Y(n18862) );
  OAI21X1 U17648 ( .A0(n25767), .A1(n26269), .B0(n17477), .Y(M4_a_20_) );
  INVX1 U17649 ( .A(n17626), .Y(n5869) );
  XNOR2X2 U17650 ( .A(n14613), .B(n14612), .Y(n20327) );
  ADDFHX2 U17651 ( .A(n17853), .B(n17852), .CI(n17851), .CO(n18410), .S(n18408) );
  AOI21X1 U17652 ( .A0(n12818), .A1(n12817), .B0(n12816), .Y(n12819) );
  ADDFX2 U17653 ( .A(n12653), .B(n12652), .CI(n12651), .CO(n12664), .S(n12679)
         );
  INVX1 U17654 ( .A(n14669), .Y(n19096) );
  NAND2X4 U17655 ( .A(n4861), .B(n4858), .Y(n14476) );
  AOI21X4 U17656 ( .A0(n13982), .A1(n14397), .B0(n5023), .Y(n4858) );
  NAND3X2 U17657 ( .A(n14578), .B(n19090), .C(n3141), .Y(n23709) );
  BUFX3 U17658 ( .A(n9838), .Y(n9974) );
  BUFX3 U17659 ( .A(n18539), .Y(n5893) );
  OAI222X1 U17660 ( .A0(n26533), .A1(n23884), .B0(n3121), .B1(n24157), .C0(
        n4582), .C1(n24616), .Y(n2599) );
  AOI21X1 U17661 ( .A0(n7808), .A1(n7807), .B0(n7806), .Y(n7809) );
  INVX8 U17662 ( .A(n20993), .Y(n19104) );
  OAI22X1 U17663 ( .A0(n18177), .A1(n18224), .B0(n18067), .B1(n18223), .Y(
        n18088) );
  OAI21X4 U17664 ( .A0(n19014), .A1(n19002), .B0(n19001), .Y(n19005) );
  XOR3X2 U17665 ( .A(n18282), .B(n18281), .C(n18280), .Y(n18283) );
  OAI21XL U17666 ( .A0(n18281), .A1(n18282), .B0(n18280), .Y(n5424) );
  INVX8 U17667 ( .A(n9050), .Y(n9164) );
  NAND2X1 U17668 ( .A(n23707), .B(n14726), .Y(n14727) );
  OAI22X1 U17669 ( .A0(n13650), .A1(n13790), .B0(n13694), .B1(n13721), .Y(
        n13688) );
  CLKINVX3 U17670 ( .A(n3214), .Y(n13605) );
  NOR2X1 U17671 ( .A(n20367), .B(n20760), .Y(n20371) );
  NOR2X1 U17672 ( .A(n4581), .B(n6229), .Y(n24266) );
  AOI21XL U17673 ( .A0(n19719), .A1(n19952), .B0(n3164), .Y(n19718) );
  XNOR2X1 U17674 ( .A(n20059), .B(n20045), .Y(n20196) );
  NOR2X1 U17675 ( .A(n19730), .B(n19807), .Y(n19662) );
  OAI21X1 U17676 ( .A0(n19358), .A1(n19361), .B0(n19359), .Y(n19401) );
  OAI21XL U17677 ( .A0(n19119), .A1(n19118), .B0(n19117), .Y(n19124) );
  OAI2BB1X2 U17678 ( .A0N(n25343), .A1N(n24064), .B0(n20168), .Y(n24070) );
  INVX1 U17679 ( .A(n25004), .Y(n25371) );
  NAND2X4 U17680 ( .A(n7885), .B(cs[2]), .Y(n21111) );
  AOI21XL U17681 ( .A0(n18298), .A1(n18297), .B0(n18296), .Y(n18311) );
  ADDFHX1 U17682 ( .A(n18279), .B(n18278), .CI(n18277), .CO(n18284), .S(n18286) );
  AOI22X2 U17683 ( .A0(n3081), .A1(n23631), .B0(n23630), .B1(n4267), .Y(n24626) );
  AOI22X2 U17684 ( .A0(n5297), .A1(n3128), .B0(n23536), .B1(n23534), .Y(n24868) );
  AOI2BB1X2 U17685 ( .A0N(n13467), .A1N(n13466), .B0(n4633), .Y(n5159) );
  OAI21X1 U17686 ( .A0(n10194), .A1(n10243), .B0(n10193), .Y(n10196) );
  AOI21X4 U17687 ( .A0(n10209), .A1(n10135), .B0(n5236), .Y(n10182) );
  AOI22XL U17688 ( .A0(n24220), .A1(n23794), .B0(temp1[15]), .B1(n2984), .Y(
        n20314) );
  NAND2X1 U17689 ( .A(n12770), .B(n12769), .Y(n12862) );
  AOI21X4 U17690 ( .A0(n10181), .A1(n5198), .B0(n5197), .Y(n10656) );
  NAND2X2 U17691 ( .A(n10480), .B(n10612), .Y(n10647) );
  OAI21XL U17692 ( .A0(n24147), .A1(n3111), .B0(n24146), .Y(n24148) );
  OAI21XL U17693 ( .A0(n24515), .A1(n3121), .B0(n23475), .Y(n2608) );
  NOR2X1 U17694 ( .A(n20929), .B(n20921), .Y(n20922) );
  OAI21X4 U17695 ( .A0(n14639), .A1(n14636), .B0(n14640), .Y(n6066) );
  OAI21X2 U17696 ( .A0(n12915), .A1(n12922), .B0(n12923), .Y(n4947) );
  OAI21XL U17697 ( .A0(n18375), .A1(n18376), .B0(n18374), .Y(n4868) );
  XOR2X1 U17698 ( .A(n18376), .B(n18375), .Y(n4871) );
  OAI222X1 U17699 ( .A0(n26525), .A1(n23884), .B0(n3121), .B1(n24226), .C0(
        n4583), .C1(n24843), .Y(n2583) );
  XOR2X2 U17700 ( .A(n5709), .B(n17472), .Y(n20939) );
  CMPR22X1 U17701 ( .A(n17680), .B(n17679), .CO(n17706), .S(n18345) );
  NAND2X1 U17702 ( .A(n4937), .B(n4936), .Y(n4935) );
  INVX4 U17703 ( .A(n9878), .Y(n9886) );
  OAI22X1 U17704 ( .A0(n9979), .A1(n9978), .B0(n9977), .B1(n9976), .Y(n9988)
         );
  NOR2X1 U17705 ( .A(n10036), .B(n10035), .Y(n10039) );
  XNOR2X2 U17706 ( .A(n14528), .B(n14527), .Y(n14686) );
  OAI22XL U17707 ( .A0(n9504), .A1(n9573), .B0(n10496), .B1(n10157), .Y(n10156) );
  XOR3X2 U17708 ( .A(n13927), .B(n13928), .C(n13926), .Y(n13923) );
  CLKINVX3 U17709 ( .A(n10718), .Y(n6142) );
  CLKINVX3 U17710 ( .A(n17483), .Y(n23736) );
  NAND2X1 U17711 ( .A(n9068), .B(n11541), .Y(M2_b_19_) );
  OAI22X1 U17712 ( .A0(n10296), .A1(n9459), .B0(n9959), .B1(n9516), .Y(n9515)
         );
  XNOR2X1 U17713 ( .A(n18503), .B(M3_mult_x_15_b_21_), .Y(n17743) );
  AOI21X1 U17714 ( .A0(n18963), .A1(n18962), .B0(n18961), .Y(n18964) );
  XOR3X2 U17715 ( .A(n5808), .B(n15999), .C(n16000), .Y(n16060) );
  XNOR2X1 U17716 ( .A(n9841), .B(n10341), .Y(n9612) );
  XOR2X2 U17717 ( .A(n5036), .B(n17599), .Y(n17691) );
  AOI21X1 U17718 ( .A0(n18318), .A1(n18317), .B0(n4668), .Y(n18327) );
  NAND2X1 U17719 ( .A(n23744), .B(n23710), .Y(n23712) );
  OAI21XL U17720 ( .A0(n12216), .A1(n12217), .B0(n4881), .Y(n4878) );
  NOR2X1 U17721 ( .A(n12851), .B(n12839), .Y(n4891) );
  NAND2XL U17722 ( .A(n21166), .B(n4722), .Y(n4894) );
  AOI21XL U17723 ( .A0(n21166), .A1(n4728), .B0(n4898), .Y(n4897) );
  AOI21XL U17724 ( .A0(n21166), .A1(n4731), .B0(n4900), .Y(n4899) );
  XNOR2X4 U17725 ( .A(M3_mult_x_15_a_17_), .B(n4918), .Y(n12746) );
  OAI2BB1X1 U17726 ( .A0N(n11835), .A1N(n4926), .B0(n4922), .Y(n11838) );
  NAND2X2 U17727 ( .A(n13986), .B(n13985), .Y(n14640) );
  NOR2X4 U17728 ( .A(n13986), .B(n13985), .Y(n14639) );
  NOR2BXL U17729 ( .AN(n24480), .B(n4935), .Y(n2458) );
  NAND2XL U17730 ( .A(n5246), .B(n25675), .Y(n4937) );
  XOR2X4 U17731 ( .A(M5_a_6_), .B(n16605), .Y(n16332) );
  XNOR2X1 U17732 ( .A(n4784), .B(n16605), .Y(n15946) );
  AOI2BB1X4 U17733 ( .A0N(n25813), .A1N(n25926), .B0(n4941), .Y(n16605) );
  XOR2X2 U17734 ( .A(M3_a_20_), .B(n12731), .Y(n11749) );
  NAND2X2 U17735 ( .A(n12501), .B(n12500), .Y(n12931) );
  NAND2X2 U17736 ( .A(n12504), .B(n12925), .Y(n12890) );
  NAND2XL U17737 ( .A(n21166), .B(n4729), .Y(n4964) );
  XOR2X2 U17738 ( .A(n12894), .B(n4629), .Y(n20321) );
  XOR2X1 U17739 ( .A(n12118), .B(n4984), .Y(n12145) );
  OAI21X1 U17740 ( .A0(n12618), .A1(n3191), .B0(n4985), .Y(n4984) );
  INVXL U17741 ( .A(n5366), .Y(n24149) );
  OAI22X1 U17742 ( .A0(n11957), .A1(n12616), .B0(n12618), .B1(n4995), .Y(
        n11944) );
  AOI21XL U17743 ( .A0(n25753), .A1(n25675), .B0(n5001), .Y(n2477) );
  XOR2X4 U17744 ( .A(n5012), .B(n20713), .Y(n20716) );
  OR2X2 U17745 ( .A(n10426), .B(n10427), .Y(n5005) );
  XOR3X2 U17746 ( .A(n10427), .B(n10425), .C(n10426), .Y(n10471) );
  NOR2X1 U17747 ( .A(n20704), .B(n20703), .Y(n20705) );
  XNOR2X4 U17748 ( .A(n5006), .B(n4681), .Y(n20614) );
  OAI2BB1X2 U17749 ( .A0N(n3132), .A1N(n20613), .B0(n20614), .Y(n5010) );
  NOR2X1 U17750 ( .A(n3078), .B(n20614), .Y(n5011) );
  NAND2X2 U17751 ( .A(n5014), .B(n4663), .Y(M4_a_18_) );
  INVXL U17752 ( .A(n17593), .Y(n5021) );
  NAND2BX1 U17753 ( .AN(n17593), .B(n3098), .Y(n5022) );
  XNOR2X4 U17754 ( .A(M1_b_22_), .B(n23173), .Y(n14356) );
  NAND2X4 U17755 ( .A(n13507), .B(n13508), .Y(n23173) );
  NAND3BX2 U17756 ( .AN(n5033), .B(n19044), .C(n23734), .Y(n5030) );
  BUFX2 U17757 ( .A(n11479), .Y(n5032) );
  OAI21XL U17758 ( .A0(n5923), .A1(n17591), .B0(n17590), .Y(n5922) );
  XOR2X1 U17759 ( .A(n17541), .B(n17540), .Y(n17590) );
  OAI22XL U17760 ( .A0(n15961), .A1(n16977), .B0(n3105), .B1(n5037), .Y(n16123) );
  XOR2X1 U17761 ( .A(n16160), .B(n16159), .Y(n5042) );
  AOI21XL U17762 ( .A0(n24655), .A1(n25754), .B0(n5043), .Y(n2319) );
  NOR2X2 U17763 ( .A(n5048), .B(n5047), .Y(n5046) );
  INVXL U17764 ( .A(n17327), .Y(n17313) );
  AOI21X4 U17765 ( .A0(n17381), .A1(n17380), .B0(n17379), .Y(n5058) );
  NAND2XL U17766 ( .A(n5061), .B(n5066), .Y(n5065) );
  NOR2X4 U17767 ( .A(n23643), .B(n5738), .Y(n25219) );
  NOR2X4 U17768 ( .A(n23643), .B(n5739), .Y(n25220) );
  OAI21XL U17769 ( .A0(n5069), .A1(n9316), .B0(n9315), .Y(n5068) );
  XOR2X2 U17770 ( .A(n5072), .B(n5071), .Y(n9414) );
  INVX1 U17771 ( .A(n9315), .Y(n5071) );
  INVX1 U17772 ( .A(n9247), .Y(n5073) );
  AOI21X4 U17773 ( .A0(n5076), .A1(n5075), .B0(n5217), .Y(n5518) );
  NAND4X2 U17774 ( .A(n5232), .B(n5231), .C(n5233), .D(n5247), .Y(n5076) );
  XOR2X4 U17775 ( .A(n5255), .B(n5079), .Y(n10329) );
  AOI22X2 U17776 ( .A0(n5297), .A1(n19104), .B0(n20615), .B1(n3128), .Y(n24913) );
  AOI22X2 U17777 ( .A0(n20712), .A1(n3128), .B0(n20615), .B1(n23722), .Y(
        n25382) );
  NOR2XL U17778 ( .A(n20686), .B(n5084), .Y(n2457) );
  AOI21XL U17779 ( .A0(n3200), .A1(n17038), .B0(n5086), .Y(
        M5_U3_U1_enc_tree_0__1__14_) );
  XOR2X4 U17780 ( .A(n16909), .B(n5086), .Y(n17061) );
  NOR2XL U17781 ( .A(n17039), .B(n5086), .Y(M5_U3_U1_enc_tree_1__1__14_) );
  OAI22X2 U17782 ( .A0(n4860), .A1(n25917), .B0(n26274), .B1(n17167), .Y(n5088) );
  NAND2X1 U17783 ( .A(target_temp[3]), .B(n9164), .Y(n5089) );
  XOR2X4 U17784 ( .A(n5091), .B(n4588), .Y(n17419) );
  XNOR3X2 U17785 ( .A(n5095), .B(n17065), .C(n17066), .Y(n17127) );
  OAI21X4 U17786 ( .A0(n26247), .A1(n25796), .B0(n5679), .Y(n17073) );
  NOR2X1 U17787 ( .A(n17133), .B(n17309), .Y(n17370) );
  AOI21X1 U17788 ( .A0(n5098), .A1(n10725), .B0(n5610), .Y(n5609) );
  INVX4 U17789 ( .A(n10727), .Y(n5098) );
  BUFX12 U17790 ( .A(n5125), .Y(n5100) );
  OAI21X4 U17791 ( .A0(n20954), .A1(n19059), .B0(n19060), .Y(n5125) );
  AOI21XL U17792 ( .A0(n24514), .A1(in_valid_d), .B0(n23730), .Y(n23731) );
  OAI2BB1X2 U17793 ( .A0N(n3455), .A1N(n20907), .B0(n5104), .Y(n24514) );
  NAND2X1 U17794 ( .A(n5604), .B(w2[5]), .Y(n5620) );
  XOR2X1 U17795 ( .A(n5105), .B(n7140), .Y(n7168) );
  OAI22XL U17796 ( .A0(n6315), .A1(n7695), .B0(n5124), .B1(n7644), .Y(n6337)
         );
  OAI22XL U17797 ( .A0(n7532), .A1(n7695), .B0(n5124), .B1(n7508), .Y(n7527)
         );
  OAI21XL U17798 ( .A0(n7546), .A1(n5124), .B0(n5107), .Y(n7566) );
  OAI22XL U17799 ( .A0(n7467), .A1(n5124), .B0(n7508), .B1(n7695), .Y(n7501)
         );
  OAI21XL U17800 ( .A0(n7532), .A1(n5124), .B0(n5108), .Y(n7551) );
  OAI22XL U17801 ( .A0(n5124), .A1(n7563), .B0(n7588), .B1(n7695), .Y(n7585)
         );
  OAI2BB2XL U17802 ( .B0(n5124), .B1(n25870), .A0N(n5122), .A1N(n25870), .Y(
        n7694) );
  NAND2BXL U17803 ( .AN(n6923), .B(n3188), .Y(n5111) );
  OAI21XL U17804 ( .A0(n7227), .A1(n5124), .B0(n5118), .Y(n7294) );
  OAI22XL U17805 ( .A0(n6824), .A1(n5124), .B0(n7695), .B1(n6842), .Y(n6838)
         );
  OAI21X1 U17806 ( .A0(n7053), .A1(n5124), .B0(n5119), .Y(n7116) );
  OAI21XL U17807 ( .A0(n6788), .A1(n5124), .B0(n5121), .Y(n6851) );
  OAI22XL U17808 ( .A0(n7695), .A1(n6784), .B0(n6346), .B1(n5124), .Y(n6759)
         );
  OAI22XL U17809 ( .A0(n7695), .A1(n6788), .B0(n6784), .B1(n5124), .Y(n6793)
         );
  NAND2X4 U17810 ( .A(n7695), .B(n6282), .Y(n5124) );
  OAI21X2 U17811 ( .A0(n7429), .A1(n7424), .B0(n7430), .Y(n7444) );
  NOR2X4 U17812 ( .A(n7264), .B(n7265), .Y(n7429) );
  NAND2X4 U17813 ( .A(n20952), .B(n20951), .Y(n20954) );
  NAND2X1 U17814 ( .A(n5128), .B(n5126), .Y(n7451) );
  OAI21X2 U17815 ( .A0(n7312), .A1(n7324), .B0(n7313), .Y(n5127) );
  OAI21X4 U17816 ( .A0(n7257), .A1(n7256), .B0(n7255), .Y(n7321) );
  OAI21X1 U17817 ( .A0(n7093), .A1(n5131), .B0(n5129), .Y(n6871) );
  NAND2X1 U17818 ( .A(n7389), .B(target_temp[18]), .Y(n5133) );
  NAND2X1 U17819 ( .A(n5135), .B(n5134), .Y(n6979) );
  NAND2XL U17820 ( .A(n5136), .B(n6951), .Y(n5135) );
  XOR2X1 U17821 ( .A(n6951), .B(n6952), .Y(n5137) );
  NAND2X2 U17822 ( .A(n5141), .B(n5140), .Y(n9688) );
  XOR2X1 U17823 ( .A(n9676), .B(n5148), .Y(n5147) );
  NAND2X2 U17824 ( .A(n14001), .B(n14595), .Y(n5280) );
  NOR2X4 U17825 ( .A(n14598), .B(n14585), .Y(n14001) );
  NOR2X4 U17826 ( .A(n13981), .B(n14399), .Y(n13982) );
  XOR3X2 U17827 ( .A(n13610), .B(n13612), .C(n13611), .Y(n13625) );
  NAND2X4 U17828 ( .A(n13972), .B(n13048), .Y(n13971) );
  XOR2X4 U17829 ( .A(n13898), .B(n5152), .Y(n13972) );
  NOR2X1 U17830 ( .A(n20999), .B(n4672), .Y(n2460) );
  XOR2X1 U17831 ( .A(n14185), .B(n5156), .Y(n14179) );
  XOR2X1 U17832 ( .A(n14187), .B(n14186), .Y(n5156) );
  NAND2X2 U17833 ( .A(n23480), .B(n23481), .Y(n23482) );
  NAND2X1 U17834 ( .A(target_temp[1]), .B(n9164), .Y(n5158) );
  NAND2XL U17835 ( .A(n13211), .B(n5164), .Y(n5160) );
  NAND2BXL U17836 ( .AN(n13211), .B(n5162), .Y(n5161) );
  XOR2X1 U17837 ( .A(n13211), .B(n5164), .Y(n5163) );
  NAND2X1 U17838 ( .A(n5165), .B(n4644), .Y(n5164) );
  NAND2X4 U17839 ( .A(n13791), .B(n5167), .Y(n13790) );
  XOR2X2 U17840 ( .A(n13605), .B(n5168), .Y(n13791) );
  OAI2BB1X2 U17841 ( .A0N(n5170), .A1N(n9518), .B0(n5169), .Y(n9528) );
  XNOR2X1 U17842 ( .A(n9519), .B(n9520), .Y(n5172) );
  NOR2XL U17843 ( .A(n5216), .B(n5175), .Y(n20945) );
  INVXL U17844 ( .A(n10703), .Y(n5175) );
  NAND2XL U17845 ( .A(n11536), .B(n4719), .Y(n5180) );
  NAND2X1 U17846 ( .A(n11536), .B(sigma10[11]), .Y(n5181) );
  XNOR2X1 U17847 ( .A(n9796), .B(n5187), .Y(n9824) );
  AOI22X2 U17848 ( .A0(y10[21]), .A1(n14427), .B0(n25229), .B1(y12[21]), .Y(
        n5189) );
  INVXL U17849 ( .A(n9649), .Y(n5196) );
  OAI21X4 U17850 ( .A0(n10182), .A1(n10144), .B0(n5234), .Y(n5197) );
  OAI21X4 U17851 ( .A0(n10278), .A1(n10127), .B0(n10126), .Y(n10181) );
  NOR2X4 U17852 ( .A(n10179), .B(n10144), .Y(n5198) );
  NAND2X1 U17853 ( .A(n11536), .B(n4727), .Y(n5200) );
  AOI22X1 U17854 ( .A0(y10[19]), .A1(n14427), .B0(n25229), .B1(y12[19]), .Y(
        n5201) );
  NAND2X4 U17855 ( .A(n9072), .B(n5203), .Y(M2_a_17_) );
  NAND2X1 U17856 ( .A(n5207), .B(n4600), .Y(n2591) );
  NAND2X1 U17857 ( .A(n20709), .B(n3132), .Y(n5209) );
  NAND2X4 U17858 ( .A(n6057), .B(n14081), .Y(n14080) );
  NAND2X1 U17859 ( .A(n5213), .B(n5212), .Y(n13759) );
  OAI21XL U17860 ( .A0(n13731), .A1(n5214), .B0(n13730), .Y(n5213) );
  AOI22X1 U17861 ( .A0(y12[13]), .A1(n4856), .B0(n14427), .B1(y10[13]), .Y(
        n5218) );
  NOR2X2 U17862 ( .A(n10320), .B(n10319), .Y(n10465) );
  NAND2X1 U17863 ( .A(n5225), .B(n5224), .Y(n10174) );
  OR2X2 U17864 ( .A(n9569), .B(n9568), .Y(n5226) );
  XOR3X2 U17865 ( .A(n9568), .B(n9569), .C(n9567), .Y(n9565) );
  NOR2X2 U17866 ( .A(n10465), .B(n10446), .Y(n10612) );
  NAND2X4 U17867 ( .A(n10190), .B(n5235), .Y(n10144) );
  NAND2XL U17868 ( .A(n9248), .B(n5245), .Y(n5241) );
  NAND2BXL U17869 ( .AN(n9248), .B(n5243), .Y(n5242) );
  INVXL U17870 ( .A(n5245), .Y(n5243) );
  XOR2X4 U17871 ( .A(n21055), .B(n5250), .Y(n10369) );
  INVX8 U17872 ( .A(n9050), .Y(n25229) );
  XNOR2X2 U17873 ( .A(n5767), .B(n3817), .Y(n23925) );
  INVXL U17874 ( .A(n10551), .Y(n10640) );
  NAND2X1 U17875 ( .A(n5260), .B(n5259), .Y(n13486) );
  CLKINVX4 U17876 ( .A(n6210), .Y(n14030) );
  NAND2X4 U17877 ( .A(target_temp[9]), .B(n4856), .Y(n13040) );
  AOI2BB1X4 U17878 ( .A0N(n14623), .A1N(n5280), .B0(n5277), .Y(n5276) );
  NAND2BX2 U17879 ( .AN(n14000), .B(n5278), .Y(n5277) );
  NAND2X1 U17880 ( .A(n6142), .B(n6141), .Y(n5281) );
  XOR2X1 U17881 ( .A(n9825), .B(n9824), .Y(n5285) );
  CLKINVX8 U17882 ( .A(n13042), .Y(n14044) );
  XNOR3X4 U17883 ( .A(n5286), .B(n13602), .C(n13604), .Y(n13685) );
  NAND2X1 U17884 ( .A(n5288), .B(n5287), .Y(n13661) );
  XOR2X1 U17885 ( .A(n5293), .B(n13751), .Y(n13817) );
  XOR2X1 U17886 ( .A(n13753), .B(n13752), .Y(n5293) );
  NAND2XL U17887 ( .A(n3066), .B(w1[135]), .Y(n5294) );
  NAND2X1 U17888 ( .A(n9164), .B(target_temp[7]), .Y(n11504) );
  OAI22X1 U17889 ( .A0(n9961), .A1(n9963), .B0(n3180), .B1(n5296), .Y(n9819)
         );
  XOR2X2 U17890 ( .A(n17488), .B(n20269), .Y(n5297) );
  XOR2XL U17891 ( .A(M2_b_15_), .B(n10540), .Y(n10336) );
  XOR2XL U17892 ( .A(n10515), .B(n10540), .Y(n10493) );
  XOR2XL U17893 ( .A(M2_mult_x_15_n1669), .B(n10540), .Y(n10512) );
  XOR2XL U17894 ( .A(n10538), .B(n10540), .Y(n10458) );
  XOR2XL U17895 ( .A(n10539), .B(n10540), .Y(n10402) );
  XOR2XL U17896 ( .A(n10335), .B(n10540), .Y(n10362) );
  XOR2XL U17897 ( .A(n10514), .B(n10540), .Y(n10379) );
  OAI21X2 U17898 ( .A0(n10541), .A1(n9360), .B0(n5305), .Y(n5304) );
  NAND2BX1 U17899 ( .AN(n9462), .B(n5758), .Y(n5305) );
  INVXL U17900 ( .A(n5306), .Y(n20807) );
  NAND2X1 U17901 ( .A(n5308), .B(n5307), .Y(n9407) );
  OAI21XL U17902 ( .A0(n9414), .A1(n9415), .B0(n9413), .Y(n5308) );
  AOI22XL U17903 ( .A0(n23794), .A1(n5312), .B0(temp1[7]), .B1(n2984), .Y(
        n20979) );
  INVXL U17904 ( .A(n5310), .Y(n2271) );
  AOI21X1 U17905 ( .A0(n25329), .A1(n5312), .B0(n24151), .Y(n5311) );
  XOR2X4 U17906 ( .A(n5314), .B(n5313), .Y(n20754) );
  NAND2X1 U17907 ( .A(n6058), .B(n19073), .Y(n5318) );
  NAND2X1 U17908 ( .A(n5322), .B(n5321), .Y(n11710) );
  NAND2XL U17909 ( .A(n11686), .B(n5964), .Y(n5321) );
  XOR2X2 U17910 ( .A(n13810), .B(n13807), .Y(n5327) );
  OAI22XL U17911 ( .A0(n16961), .A1(n16960), .B0(n16962), .B1(n5329), .Y(
        n16958) );
  NOR2X4 U17912 ( .A(n14603), .B(n14609), .Y(n14595) );
  NAND2X1 U17913 ( .A(n13596), .B(n13595), .Y(n14400) );
  NOR2X4 U17914 ( .A(n13646), .B(n13645), .Y(n13981) );
  INVX1 U17915 ( .A(n16301), .Y(n5333) );
  XOR2X2 U17916 ( .A(n20689), .B(n20688), .Y(n23882) );
  XOR2X4 U17917 ( .A(n14729), .B(n4752), .Y(n20690) );
  NAND2X1 U17918 ( .A(n25229), .B(y12[5]), .Y(n5347) );
  OAI21XL U17919 ( .A0(n9285), .A1(n9284), .B0(n9283), .Y(n5350) );
  NOR2X2 U17920 ( .A(n7447), .B(n7438), .Y(n5354) );
  NAND2X1 U17921 ( .A(n5360), .B(n5359), .Y(n7196) );
  OAI21XL U17922 ( .A0(n7219), .A1(n7460), .B0(n5361), .Y(n7225) );
  NAND2XL U17923 ( .A(n5363), .B(n5362), .Y(n5361) );
  XOR2X1 U17924 ( .A(n23220), .B(n25875), .Y(n5363) );
  NAND2XL U17925 ( .A(n11977), .B(n5373), .Y(n5368) );
  NAND2XL U17926 ( .A(n5370), .B(n11976), .Y(n5369) );
  INVXL U17927 ( .A(n5373), .Y(n5371) );
  NAND2X1 U17928 ( .A(n3008), .B(n5380), .Y(n5379) );
  NAND2X1 U17929 ( .A(n23743), .B(n5388), .Y(n5382) );
  NAND2BX1 U17930 ( .AN(n23743), .B(n5384), .Y(n5383) );
  NOR2X2 U17931 ( .A(n5396), .B(n7768), .Y(n7668) );
  XOR2X2 U17932 ( .A(n25869), .B(n5398), .Y(n6292) );
  XNOR2X1 U17933 ( .A(n12442), .B(n12444), .Y(n5405) );
  NAND2X1 U17934 ( .A(n5408), .B(n25807), .Y(n5407) );
  NAND2X4 U17935 ( .A(n4674), .B(n5411), .Y(M3_mult_x_15_b_20_) );
  NAND2XL U17936 ( .A(n5413), .B(n12631), .Y(n5412) );
  OAI21X4 U17937 ( .A0(n4860), .A1(n25910), .B0(n5417), .Y(M3_mult_x_15_a_17_)
         );
  INVXL U17938 ( .A(n18292), .Y(n5421) );
  NOR2X1 U17939 ( .A(n18293), .B(n18292), .Y(n18295) );
  NOR2X1 U17940 ( .A(n5429), .B(n3015), .Y(n5426) );
  NAND2X4 U17941 ( .A(n5432), .B(n5431), .Y(M3_mult_x_15_n1682) );
  XNOR2X1 U17942 ( .A(n3022), .B(n5430), .Y(n16203) );
  XNOR2X1 U17943 ( .A(n18550), .B(n5444), .Y(n5443) );
  AOI2BB1X2 U17944 ( .A0N(n18434), .A1N(n3195), .B0(n5445), .Y(n5444) );
  OR2X2 U17945 ( .A(n17907), .B(n18107), .Y(n5447) );
  OR2XL U17946 ( .A(n17906), .B(n18235), .Y(n5448) );
  NAND2BX1 U17947 ( .AN(n5452), .B(n20700), .Y(n5451) );
  INVX1 U17948 ( .A(n23549), .Y(n5454) );
  XOR2X1 U17949 ( .A(n5430), .B(n18106), .Y(n5460) );
  NOR2X1 U17950 ( .A(n18211), .B(n18210), .Y(n5461) );
  OAI21X2 U17951 ( .A0(n5769), .A1(n18541), .B0(n5768), .Y(n17720) );
  MXI2X4 U17952 ( .A(n5462), .B(M4_a_12_), .S0(n18428), .Y(n18539) );
  OAI22X1 U17953 ( .A0(n18223), .A1(n5466), .B0(n18112), .B1(n18177), .Y(
        n18115) );
  AOI22X2 U17954 ( .A0(n3128), .A1(n5478), .B0(n23462), .B1(n23534), .Y(n24536) );
  OAI21X4 U17955 ( .A0(n25767), .A1(n26252), .B0(n5481), .Y(M4_a_13_) );
  XOR2X4 U17956 ( .A(n5484), .B(n14548), .Y(n20665) );
  XOR2X4 U17957 ( .A(n5485), .B(n14540), .Y(n14689) );
  NAND2X2 U17958 ( .A(target_temp[13]), .B(n25229), .Y(n5504) );
  XOR3X2 U17959 ( .A(n14056), .B(n14054), .C(n14055), .Y(n14068) );
  CLKINVX2 U17960 ( .A(n14532), .Y(n5501) );
  NOR2X1 U17961 ( .A(n5507), .B(n18625), .Y(n6084) );
  XOR2X1 U17962 ( .A(M3_mult_x_15_n1682), .B(n18603), .Y(n5507) );
  OAI22X1 U17963 ( .A0(n18083), .A1(n4649), .B0(n18429), .B1(n17870), .Y(
        n17891) );
  NOR2X4 U17964 ( .A(n5511), .B(n5513), .Y(n14119) );
  NAND2XL U17965 ( .A(n21166), .B(sigma11[23]), .Y(n18739) );
  NAND2XL U17966 ( .A(n21166), .B(sigma11[24]), .Y(n18741) );
  NAND2XL U17967 ( .A(n21166), .B(sigma12[23]), .Y(n17157) );
  NAND2XL U17968 ( .A(n21166), .B(sigma12[24]), .Y(n17160) );
  NAND2XL U17969 ( .A(n21166), .B(sigma11[26]), .Y(n18747) );
  NAND2XL U17970 ( .A(n21166), .B(sigma12[26]), .Y(n17166) );
  NAND2XL U17971 ( .A(n21166), .B(sigma12[28]), .Y(n17173) );
  NAND2XL U17972 ( .A(n21166), .B(sigma12[30]), .Y(n17154) );
  NAND2XL U17973 ( .A(n21166), .B(sigma11[25]), .Y(n18745) );
  NAND2XL U17974 ( .A(n21166), .B(target_temp[24]), .Y(n11598) );
  NAND2XL U17975 ( .A(n21166), .B(target_temp[23]), .Y(n11601) );
  NAND2XL U17976 ( .A(n21166), .B(sigma12[25]), .Y(n17164) );
  NAND2XL U17977 ( .A(n21166), .B(sigma11[27]), .Y(n18751) );
  NAND2XL U17978 ( .A(n21166), .B(sigma12[27]), .Y(n17171) );
  NAND2XL U17979 ( .A(n21166), .B(sigma12[29]), .Y(n17177) );
  NAND2XL U17980 ( .A(n21166), .B(sigma11[31]), .Y(n22479) );
  NAND2X1 U17981 ( .A(n5514), .B(n24215), .Y(n24216) );
  AND2X2 U17982 ( .A(n23557), .B(n23734), .Y(n5515) );
  NAND2X1 U17983 ( .A(n14317), .B(n14318), .Y(n14563) );
  XOR2X1 U17984 ( .A(n9841), .B(M2_b_15_), .Y(n5517) );
  OAI21X2 U17985 ( .A0(n5522), .A1(n5521), .B0(n5520), .Y(n9527) );
  XOR2X2 U17986 ( .A(n5525), .B(n5524), .Y(n5523) );
  NAND2X2 U17987 ( .A(n10125), .B(n10197), .Y(n10127) );
  XOR2X1 U17988 ( .A(n10290), .B(n10291), .Y(n5529) );
  XOR2X1 U17989 ( .A(n9422), .B(n5534), .Y(n5530) );
  NAND2XL U17990 ( .A(n9423), .B(n5534), .Y(n5531) );
  INVXL U17991 ( .A(n9445), .Y(n5538) );
  XOR2X4 U17992 ( .A(n10322), .B(n4626), .Y(n17482) );
  OAI21XL U17993 ( .A0(n5859), .A1(n5545), .B0(n16411), .Y(n5856) );
  OAI21XL U17994 ( .A0(n24352), .A1(n3121), .B0(n5560), .Y(n2566) );
  NOR2X4 U17995 ( .A(n7004), .B(n7003), .Y(n7257) );
  NOR2X4 U17996 ( .A(n7261), .B(n7260), .Y(n7312) );
  NAND2X1 U17997 ( .A(n7266), .B(n7267), .Y(n7448) );
  NAND2X4 U17998 ( .A(n7556), .B(n5572), .Y(n7535) );
  NOR2X1 U17999 ( .A(n6266), .B(n26255), .Y(n5581) );
  NAND2BX4 U18000 ( .AN(n5583), .B(n5627), .Y(n6613) );
  NAND3BX1 U18001 ( .AN(n20364), .B(n20366), .C(n5585), .Y(n20367) );
  OAI22X4 U18002 ( .A0(n5590), .A1(n5589), .B0(n5587), .B1(n5586), .Y(n25828)
         );
  XOR2X2 U18003 ( .A(n5592), .B(n5591), .Y(n5590) );
  NAND2X2 U18004 ( .A(n7258), .B(n7259), .Y(n7324) );
  OR2X2 U18005 ( .A(n6713), .B(n6712), .Y(n5616) );
  XOR3X2 U18006 ( .A(n6532), .B(n6533), .C(n6531), .Y(n6546) );
  NOR2X1 U18007 ( .A(n6715), .B(n6714), .Y(n6717) );
  XOR2X1 U18008 ( .A(n5634), .B(n6499), .Y(n5633) );
  NOR2X2 U18009 ( .A(n18975), .B(n18976), .Y(n5637) );
  OAI22XL U18010 ( .A0(n18483), .A1(n17636), .B0(n3195), .B1(n17734), .Y(
        n17733) );
  INVX1 U18011 ( .A(n19022), .Y(n23549) );
  OAI21X2 U18012 ( .A0(n7382), .A1(n26014), .B0(n6268), .Y(M0_a_16_) );
  XNOR2X2 U18013 ( .A(M0_a_15_), .B(M0_a_16_), .Y(n6300) );
  NOR2X1 U18014 ( .A(n17315), .B(n17316), .Y(n17311) );
  AOI22X2 U18015 ( .A0(n19104), .A1(n20754), .B0(n20814), .B1(n3128), .Y(
        n24769) );
  OAI22X1 U18016 ( .A0(n10660), .A1(n9960), .B0(n3178), .B1(n3182), .Y(n9250)
         );
  CMPR22X1 U18017 ( .A(n9251), .B(n9250), .CO(n9299), .S(n9306) );
  AOI22X1 U18018 ( .A0(n3139), .A1(n20872), .B0(n20900), .B1(n3455), .Y(n23912) );
  ADDFHX4 U18019 ( .A(n12674), .B(n12673), .CI(n12672), .CO(n12764), .S(n12511) );
  OAI22X1 U18020 ( .A0(n18541), .A1(n17510), .B0(n5893), .B1(n17623), .Y(
        n17641) );
  OAI22X1 U18021 ( .A0(n18226), .A1(n17994), .B0(n17963), .B1(n17962), .Y(
        n17993) );
  MXI2X1 U18022 ( .A(mul5_out[17]), .B(n5849), .S0(n4772), .Y(n2330) );
  OAI21X1 U18023 ( .A0(n16922), .A1(n17092), .B0(n5825), .Y(n17042) );
  XNOR2X1 U18024 ( .A(n18453), .B(M3_mult_x_15_b_9_), .Y(n17655) );
  NAND2XL U18025 ( .A(n18300), .B(n18299), .Y(n18304) );
  XOR3X2 U18026 ( .A(n17919), .B(n5811), .C(n17918), .Y(n17959) );
  AOI22XL U18027 ( .A0(n25770), .A1(n25807), .B0(n2984), .B1(temp1[29]), .Y(
        n24052) );
  AOI22XL U18028 ( .A0(n25679), .A1(n25807), .B0(n2983), .B1(temp1[26]), .Y(
        n25680) );
  NOR2X2 U18029 ( .A(n23648), .B(n20305), .Y(n20666) );
  OAI21XL U18030 ( .A0(n16758), .A1(n16757), .B0(n16756), .Y(n16759) );
  NAND2X1 U18031 ( .A(n18302), .B(n18301), .Y(n18303) );
  XOR3X2 U18032 ( .A(n18077), .B(n18076), .C(n18075), .Y(n18300) );
  OAI22XL U18033 ( .A0(n18111), .A1(n18066), .B0(n18504), .B1(n18026), .Y(
        n18065) );
  AOI21X1 U18034 ( .A0(n18896), .A1(n18900), .B0(n18887), .Y(n18888) );
  OAI21X1 U18035 ( .A0(n18889), .A1(n18925), .B0(n18888), .Y(n18894) );
  XOR2X1 U18036 ( .A(n18991), .B(n4696), .Y(n20698) );
  INVX1 U18037 ( .A(n20691), .Y(n17462) );
  XNOR2X1 U18038 ( .A(n3204), .B(n16884), .Y(n12022) );
  OAI21X2 U18039 ( .A0(n5657), .A1(n16772), .B0(n16771), .Y(n5656) );
  XNOR2X1 U18040 ( .A(n18118), .B(n3021), .Y(n17603) );
  XNOR2X2 U18041 ( .A(n3211), .B(n5645), .Y(n15944) );
  XNOR3X2 U18042 ( .A(n16303), .B(n5690), .C(n16302), .Y(n16296) );
  NAND2X1 U18043 ( .A(n16864), .B(n16865), .Y(n17246) );
  XOR2X4 U18044 ( .A(n5659), .B(n4595), .Y(n20348) );
  NAND2BXL U18045 ( .AN(n16972), .B(n5670), .Y(n5669) );
  OAI21X1 U18046 ( .A0(n16311), .A1(n17060), .B0(n5673), .Y(n5672) );
  OAI22X1 U18047 ( .A0(n16960), .A1(n3211), .B0(n16962), .B1(n5692), .Y(n16911) );
  OAI21X1 U18048 ( .A0(mul5_out[22]), .A1(n5032), .B0(n25764), .Y(n2340) );
  AOI22XL U18049 ( .A0(n5720), .A1(n17439), .B0(n17448), .B1(n5335), .Y(n17440) );
  OAI2BB1X2 U18050 ( .A0N(n16393), .A1N(n5703), .B0(n5702), .Y(n16432) );
  XOR2X2 U18051 ( .A(n5708), .B(n17423), .Y(n17430) );
  AOI21X1 U18052 ( .A0(n17210), .A1(n17211), .B0(n5713), .Y(n5712) );
  NAND2X2 U18053 ( .A(n5715), .B(n5717), .Y(n17434) );
  NOR2X4 U18054 ( .A(n5714), .B(n17420), .Y(n5715) );
  NAND4X4 U18055 ( .A(n5715), .B(n5717), .C(n5716), .D(n17433), .Y(n20929) );
  NOR2X4 U18056 ( .A(n17432), .B(n17431), .Y(n5716) );
  NOR2X1 U18057 ( .A(n17420), .B(n20340), .Y(n20735) );
  XNOR2X1 U18058 ( .A(M5_a_8_), .B(n5729), .Y(n15967) );
  INVXL U18059 ( .A(n16734), .Y(n5736) );
  NOR2BX1 U18060 ( .AN(n9722), .B(n5746), .Y(n9727) );
  NOR2X1 U18061 ( .A(n5748), .B(n5747), .Y(n5746) );
  NOR2XL U18062 ( .A(n9693), .B(n3180), .Y(n5747) );
  XOR2X1 U18063 ( .A(n20347), .B(n5750), .Y(n21048) );
  OAI22XL U18064 ( .A0(n10336), .A1(n10541), .B0(n10362), .B1(n3174), .Y(
        n10360) );
  OAI22XL U18065 ( .A0(n10541), .A1(n10493), .B0(n10512), .B1(n3174), .Y(
        n10511) );
  OAI21XL U18066 ( .A0(n10458), .A1(n10541), .B0(n5753), .Y(n10489) );
  OAI21XL U18067 ( .A0(n10541), .A1(n10512), .B0(n5754), .Y(n10530) );
  OAI21XL U18068 ( .A0(n25885), .A1(n3174), .B0(n5755), .Y(n10544) );
  OAI21XL U18069 ( .A0(n10379), .A1(n3174), .B0(n5756), .Y(n10383) );
  BUFX2 U18070 ( .A(n20698), .Y(n5771) );
  XOR2X4 U18071 ( .A(n19005), .B(n4688), .Y(n20697) );
  XOR2X2 U18072 ( .A(n5781), .B(n5780), .Y(n12041) );
  NAND2XL U18073 ( .A(n17730), .B(n5794), .Y(n5793) );
  NOR2X1 U18074 ( .A(n17620), .B(n18107), .Y(n5798) );
  NAND3X1 U18075 ( .A(n17419), .B(n5800), .C(n24259), .Y(n17235) );
  NAND2X1 U18076 ( .A(n5800), .B(n20744), .Y(n20340) );
  CLKINVX3 U18077 ( .A(n20692), .Y(n5800) );
  NAND2BXL U18078 ( .AN(n16428), .B(n5805), .Y(n5804) );
  OAI22X1 U18079 ( .A0(n16941), .A1(n16010), .B0(n15973), .B1(n16939), .Y(
        n5808) );
  OAI21X1 U18080 ( .A0(n5818), .A1(n5817), .B0(n5816), .Y(n17984) );
  INVX1 U18081 ( .A(n17971), .Y(n5817) );
  NAND2X1 U18082 ( .A(n23734), .B(n6024), .Y(n5822) );
  XNOR2X1 U18083 ( .A(n18589), .B(n18590), .Y(n5823) );
  OAI21XL U18084 ( .A0(n16922), .A1(n17099), .B0(n5826), .Y(n16921) );
  OR2XL U18085 ( .A(n16903), .B(n17092), .Y(n5826) );
  OAI21XL U18086 ( .A0(n16871), .A1(n17092), .B0(n5828), .Y(n16887) );
  OR2XL U18087 ( .A(n16889), .B(n17099), .Y(n5828) );
  NAND2X1 U18088 ( .A(n5833), .B(n5832), .Y(mul5_out[11]) );
  NOR2XL U18089 ( .A(n5835), .B(n3207), .Y(n16623) );
  OAI21XL U18090 ( .A0(n16631), .A1(n16704), .B0(n5836), .Y(n16633) );
  OAI21XL U18091 ( .A0(n16573), .A1(n5835), .B0(n5837), .Y(n16587) );
  NAND2BXL U18092 ( .AN(n16581), .B(n5847), .Y(n5837) );
  OAI21XL U18093 ( .A0(n16581), .A1(n5835), .B0(n5838), .Y(n16597) );
  OAI21XL U18094 ( .A0(n16613), .A1(n5835), .B0(n5839), .Y(n16650) );
  OAI21XL U18095 ( .A0(n16602), .A1(n5835), .B0(n5840), .Y(n16612) );
  OAI22XL U18096 ( .A0(n16381), .A1(n5835), .B0(n16343), .B1(n16704), .Y(
        n16364) );
  OAI21XL U18097 ( .A0(n16703), .A1(n5835), .B0(n5841), .Y(n16713) );
  OAI22XL U18098 ( .A0(n16640), .A1(n16704), .B0(n16639), .B1(n5835), .Y(
        n16651) );
  OAI21XL U18099 ( .A0(n16702), .A1(n5835), .B0(n5843), .Y(n16708) );
  OAI21XL U18100 ( .A0(n16702), .A1(n16704), .B0(n5844), .Y(n16705) );
  OAI21XL U18101 ( .A0(n16469), .A1(n5835), .B0(n5846), .Y(n16499) );
  NAND2X1 U18102 ( .A(n20943), .B(n5336), .Y(n5852) );
  OAI21X4 U18103 ( .A0(n5855), .A1(n5854), .B0(n5853), .Y(n16451) );
  INVX1 U18104 ( .A(n16417), .Y(n5854) );
  XOR2X1 U18105 ( .A(n16411), .B(n5859), .Y(n5858) );
  NAND2X1 U18106 ( .A(n17626), .B(n17627), .Y(n5867) );
  NAND2X1 U18107 ( .A(n5869), .B(n5870), .Y(n5868) );
  NAND2X4 U18108 ( .A(n5871), .B(n18539), .Y(n18541) );
  OAI22X1 U18109 ( .A0(n18111), .A1(n17602), .B0(n17538), .B1(n18504), .Y(
        n17591) );
  NOR2X4 U18110 ( .A(n19043), .B(n3111), .Y(n24117) );
  AND2X2 U18111 ( .A(n19049), .B(n23734), .Y(n5880) );
  OAI22X2 U18112 ( .A0(n18107), .A1(n17735), .B0(n18235), .B1(n18118), .Y(
        n5887) );
  XOR2X1 U18113 ( .A(n18943), .B(n4639), .Y(n19022) );
  XOR2X1 U18114 ( .A(n18998), .B(n4704), .Y(n23551) );
  XOR2X1 U18115 ( .A(n5904), .B(n17843), .Y(n17853) );
  XOR2X1 U18116 ( .A(n17842), .B(n17844), .Y(n5904) );
  XNOR2X1 U18117 ( .A(n17566), .B(n5909), .Y(n5908) );
  NOR2X1 U18118 ( .A(n18107), .B(n17505), .Y(n5910) );
  NAND2X1 U18119 ( .A(n23734), .B(n23477), .Y(n5921) );
  AOI21XL U18120 ( .A0(n25754), .A1(n24842), .B0(n5925), .Y(n2331) );
  NAND2X1 U18121 ( .A(n12512), .B(n12511), .Y(n12923) );
  INVXL U18122 ( .A(n5939), .Y(n5937) );
  XOR2X1 U18123 ( .A(n5938), .B(n11987), .Y(n11989) );
  XOR2X1 U18124 ( .A(n11988), .B(n5939), .Y(n5938) );
  INVXL U18125 ( .A(n20671), .Y(n20309) );
  OAI22X1 U18126 ( .A0(n12618), .A1(n5956), .B0(n12616), .B1(n25884), .Y(
        n12563) );
  INVXL U18127 ( .A(n5964), .Y(n5962) );
  XOR2X2 U18128 ( .A(n11686), .B(n5963), .Y(n11738) );
  NOR2X2 U18129 ( .A(n12897), .B(n12896), .Y(n12925) );
  XOR2X1 U18130 ( .A(n11875), .B(n11874), .Y(n5975) );
  XOR2X2 U18131 ( .A(M3_a_20_), .B(n12758), .Y(n5984) );
  NAND2X1 U18132 ( .A(n4875), .B(data[39]), .Y(n5988) );
  INVX1 U18133 ( .A(n5990), .Y(n20844) );
  XOR2X1 U18134 ( .A(n12698), .B(n5996), .Y(n5995) );
  OAI22X1 U18135 ( .A0(n12576), .A1(n12575), .B0(n12760), .B1(n12700), .Y(
        n5996) );
  NAND2BX4 U18136 ( .AN(n6156), .B(n6023), .Y(M3_mult_x_15_b_2_) );
  OAI2BB1X2 U18137 ( .A0N(n20899), .A1N(n3455), .B0(n6025), .Y(n24644) );
  XOR2X1 U18138 ( .A(M3_mult_x_15_b_1_), .B(n18428), .Y(n6026) );
  NAND2X4 U18139 ( .A(n6300), .B(n6027), .Y(n7633) );
  OAI21XL U18140 ( .A0(n18119), .A1(n18107), .B0(n6037), .Y(n18132) );
  NAND2XL U18141 ( .A(n6039), .B(n6038), .Y(n6037) );
  OR2X2 U18142 ( .A(n18201), .B(n18200), .Y(n18204) );
  NOR2XL U18143 ( .A(n17486), .B(n20810), .Y(n17487) );
  NOR2XL U18144 ( .A(M2_mult_x_15_n1669), .B(n10515), .Y(
        M2_U4_U1_enc_tree_1__1__10_) );
  AOI21XL U18145 ( .A0(M2_U4_U1_or2_inv_0__10_), .A1(M2_mult_x_15_n1668), .B0(
        n10515), .Y(M2_U4_U1_enc_tree_0__1__10_) );
  NAND2X2 U18146 ( .A(n11543), .B(n9063), .Y(n10515) );
  NAND2X4 U18147 ( .A(n6049), .B(n9049), .Y(n10341) );
  XOR2X1 U18148 ( .A(n5489), .B(n14236), .Y(n13695) );
  XNOR2X1 U18149 ( .A(n5489), .B(M1_b_10_), .Y(n6057) );
  OAI22X1 U18150 ( .A0(n9550), .A1(n9966), .B0(n10159), .B1(n9841), .Y(n9584)
         );
  NAND2X4 U18151 ( .A(n9214), .B(n10159), .Y(n9966) );
  NAND2X4 U18152 ( .A(n4580), .B(n6161), .Y(n9050) );
  XOR3X2 U18153 ( .A(n9692), .B(n9691), .C(n9690), .Y(n9764) );
  NAND2XL U18154 ( .A(n14208), .B(n14198), .Y(n6069) );
  XOR2X4 U18155 ( .A(n6070), .B(n4616), .Y(n6074) );
  NOR2X2 U18156 ( .A(n10278), .B(n10199), .Y(n6071) );
  NOR2X2 U18157 ( .A(n14690), .B(n14691), .Y(n6073) );
  XNOR2X1 U18158 ( .A(n6082), .B(n17550), .Y(n6081) );
  NOR2X1 U18159 ( .A(n18923), .B(n18919), .Y(n18903) );
  NAND2X4 U18160 ( .A(n12523), .B(n11633), .Y(n12597) );
  XOR3X2 U18161 ( .A(n14022), .B(n14021), .C(n14020), .Y(n14009) );
  OAI22X1 U18162 ( .A0(n6101), .A1(n12597), .B0(n12595), .B1(n12072), .Y(
        n12109) );
  NOR2X2 U18163 ( .A(n14309), .B(n14310), .Y(n14590) );
  NAND2X2 U18164 ( .A(n12491), .B(n12490), .Y(n12937) );
  OAI2BB1X4 U18165 ( .A0N(n6117), .A1N(n16076), .B0(n6116), .Y(n16153) );
  OAI2BB1X1 U18166 ( .A0N(n15978), .A1N(n15977), .B0(n6120), .Y(n16019) );
  OAI21XL U18167 ( .A0(n15977), .A1(n15978), .B0(n15976), .Y(n6120) );
  XNOR3X2 U18168 ( .A(n15978), .B(n15977), .C(n6121), .Y(n16058) );
  NAND2X1 U18169 ( .A(n20657), .B(n22482), .Y(n6133) );
  NAND2X1 U18170 ( .A(n6136), .B(n6135), .Y(n12383) );
  CLKINVX3 U18171 ( .A(n13720), .Y(n13693) );
  OAI22X1 U18172 ( .A0(n12152), .A1(n6137), .B0(n3185), .B1(n12353), .Y(n12362) );
  XOR2X4 U18173 ( .A(n10388), .B(M2_a_16_), .Y(n10496) );
  XOR2X1 U18174 ( .A(n16614), .B(n6146), .Y(n6145) );
  OAI21X4 U18175 ( .A0(n10283), .A1(n10280), .B0(n10284), .Y(n10198) );
  NAND2X1 U18176 ( .A(n6151), .B(n6150), .Y(n16095) );
  OAI21XL U18177 ( .A0(n4780), .A1(n16099), .B0(n16098), .Y(n6151) );
  XOR3X2 U18178 ( .A(n4780), .B(n16098), .C(n16099), .Y(n16811) );
  XOR2X1 U18179 ( .A(n10428), .B(n10430), .Y(n6165) );
  XNOR2X1 U18180 ( .A(M0_b_9_), .B(n25866), .Y(n6491) );
  AOI21X1 U18181 ( .A0(n7436), .A1(n7426), .B0(n7425), .Y(n7427) );
  ADDFHX4 U18182 ( .A(n7251), .B(n7250), .CI(n7249), .CO(n7260), .S(n7258) );
  ADDFHX1 U18183 ( .A(n6880), .B(n6879), .CI(n6878), .CO(n6953), .S(n6890) );
  CMPR22X1 U18184 ( .A(n12036), .B(n12035), .CO(n12056), .S(n12077) );
  AOI21XL U18185 ( .A0(n20268), .A1(n3060), .B0(n20267), .Y(n2468) );
  XNOR2X1 U18186 ( .A(n4567), .B(n25862), .Y(n13653) );
  OAI22X1 U18187 ( .A0(n13914), .A1(n14198), .B0(n13875), .B1(n14208), .Y(
        n13930) );
  XNOR2X1 U18188 ( .A(n25884), .B(n3021), .Y(n11957) );
  OAI21XL U18189 ( .A0(n24536), .A1(n3024), .B0(n24533), .Y(n24534) );
  OAI21XL U18190 ( .A0(n24536), .A1(n3121), .B0(n23891), .Y(n2606) );
  NAND2X2 U18191 ( .A(n11509), .B(n11508), .Y(M1_b_4_) );
  CLKINVX3 U18192 ( .A(n13057), .Y(n13843) );
  CMPR22X1 U18193 ( .A(n13551), .B(n13550), .CO(n13635), .S(n13579) );
  OAI22X1 U18194 ( .A0(n13555), .A1(n14268), .B0(n13512), .B1(n14282), .Y(
        n13550) );
  OAI21XL U18195 ( .A0(n25506), .A1(n3121), .B0(n23954), .Y(n2596) );
  INVX1 U18196 ( .A(n23912), .Y(n23658) );
  OAI22X1 U18197 ( .A0(n6988), .A1(n7633), .B0(n7026), .B1(n7634), .Y(n7072)
         );
  ADDFX2 U18198 ( .A(n11733), .B(n11732), .CI(n11731), .CO(n11741), .S(n11805)
         );
  XNOR2X1 U18199 ( .A(n3204), .B(n12803), .Y(n11914) );
  OAI22XL U18200 ( .A0(n13399), .A1(n13790), .B0(n13450), .B1(n13721), .Y(
        n13445) );
  AOI22XL U18201 ( .A0(n24350), .A1(n25807), .B0(n2984), .B1(temp2[25]), .Y(
        n24351) );
  OAI21XL U18202 ( .A0(n24352), .A1(n4582), .B0(n24351), .Y(n2567) );
  OAI22X1 U18203 ( .A0(n3102), .A1(n15964), .B0(n16332), .B1(n15959), .Y(
        n15989) );
  INVX8 U18204 ( .A(in_valid_t), .Y(n15940) );
  AOI21X1 U18205 ( .A0(n7389), .A1(y10[7]), .B0(n25145), .Y(n6247) );
  XNOR2XL U18206 ( .A(n18118), .B(n11499), .Y(n18234) );
  XNOR2X1 U18207 ( .A(n17039), .B(n3196), .Y(n16876) );
  OAI22X1 U18208 ( .A0(n6330), .A1(n7633), .B0(n6349), .B1(n7634), .Y(n6354)
         );
  OAI22X1 U18209 ( .A0(n6330), .A1(n7634), .B0(n7633), .B1(n6325), .Y(n6382)
         );
  OAI22XL U18210 ( .A0(n6988), .A1(n7634), .B0(n7633), .B1(n6941), .Y(n6987)
         );
  AOI2BB1X1 U18211 ( .A0N(n20914), .A1N(n4581), .B0(n19087), .Y(n19088) );
  XNOR2X1 U18212 ( .A(n12265), .B(n12560), .Y(n12012) );
  ADDFHX1 U18213 ( .A(n18531), .B(n18530), .CI(n18529), .CO(n18567), .S(n18571) );
  ADDFHX1 U18214 ( .A(n13546), .B(n13545), .CI(n13544), .CO(n13584), .S(n13549) );
  XOR2X1 U18215 ( .A(n10742), .B(n20276), .Y(n20882) );
  XOR2X2 U18216 ( .A(n20753), .B(n20752), .Y(n20814) );
  XNOR2X1 U18217 ( .A(n18006), .B(M3_mult_x_15_b_9_), .Y(n18225) );
  XNOR2X2 U18218 ( .A(n7751), .B(n7750), .Y(n20283) );
  AOI22XL U18219 ( .A0(n9164), .A1(y12[2]), .B0(n14427), .B1(y10[2]), .Y(n9052) );
  XNOR2X1 U18220 ( .A(n12594), .B(M3_mult_x_15_b_1_), .Y(n12201) );
  ADDFHX1 U18221 ( .A(n13853), .B(n13852), .CI(n13851), .CO(n13904), .S(n13833) );
  OAI22X1 U18222 ( .A0(n12715), .A1(n11783), .B0(n12525), .B1(n11880), .Y(
        n11890) );
  XNOR2X1 U18223 ( .A(n12732), .B(n16884), .Y(n11880) );
  AOI21X1 U18224 ( .A0(n18855), .A1(n18851), .B0(n18682), .Y(n18927) );
  ADDFHX4 U18225 ( .A(n13802), .B(n13801), .CI(n13800), .CO(n13989), .S(n13988) );
  XNOR2X1 U18226 ( .A(n3209), .B(n7800), .Y(n6963) );
  XNOR2X1 U18227 ( .A(n25883), .B(M3_mult_x_15_b_1_), .Y(n17672) );
  OAI22X1 U18228 ( .A0(n18659), .A1(n17553), .B0(n17832), .B1(n17511), .Y(
        n17498) );
  ADDFHX4 U18229 ( .A(n16266), .B(n16265), .CI(n16264), .CO(n16297), .S(n16293) );
  ADDFHX4 U18230 ( .A(n17856), .B(n17855), .CI(n17854), .CO(n18413), .S(n18411) );
  OAI22X1 U18231 ( .A0(n10368), .A1(n9381), .B0(n9780), .B1(n9252), .Y(n9377)
         );
  OAI22X1 U18232 ( .A0(n10368), .A1(n9382), .B0(n9780), .B1(n9381), .Y(n9423)
         );
  AOI22X1 U18233 ( .A0(n3139), .A1(n20819), .B0(n20847), .B1(n23892), .Y(
        n24783) );
  AOI22X1 U18234 ( .A0(n3139), .A1(n20956), .B0(n23892), .B1(n20955), .Y(
        n25687) );
  AOI22X1 U18235 ( .A0(n20907), .A1(n3139), .B0(n19079), .B1(n3455), .Y(n20914) );
  INVX4 U18236 ( .A(n13045), .Y(n13721) );
  OAI22XL U18237 ( .A0(n18111), .A1(n18227), .B0(n18504), .B1(n18086), .Y(
        n18218) );
  XNOR2X1 U18238 ( .A(n18503), .B(M3_mult_x_15_b_3_), .Y(n18086) );
  INVX4 U18239 ( .A(n10181), .Y(n10243) );
  OAI22X1 U18240 ( .A0(n18666), .A1(n18658), .B0(n17832), .B1(n17606), .Y(
        n17679) );
  ADDFHX1 U18241 ( .A(n13633), .B(n13632), .CI(n13631), .CO(n13709), .S(n13640) );
  OAI22X1 U18242 ( .A0(n17092), .A1(n16135), .B0(n16317), .B1(n16184), .Y(
        n16181) );
  XNOR2X1 U18243 ( .A(n7286), .B(n7646), .Y(n6976) );
  ADDFHX1 U18244 ( .A(n10022), .B(n10021), .CI(n10020), .CO(n10027), .S(n10029) );
  OAI21X2 U18245 ( .A0(n7382), .A1(n26013), .B0(n6259), .Y(M0_a_15_) );
  ADDFHX1 U18246 ( .A(n16234), .B(n16233), .CI(n16232), .CO(n16262), .S(n16258) );
  OAI22X1 U18247 ( .A0(n9504), .A1(n9434), .B0(n10496), .B1(n9419), .Y(n9438)
         );
  XNOR2X1 U18248 ( .A(n3209), .B(n25872), .Y(n7027) );
  ADDFHX4 U18249 ( .A(n9491), .B(n9490), .CI(n9489), .CO(n10139), .S(n10137)
         );
  AOI22X1 U18250 ( .A0(n5336), .A1(n24263), .B0(n3136), .B1(n6221), .Y(n24264)
         );
  OAI21X1 U18251 ( .A0(n3494), .A1(n7753), .B0(n7757), .Y(n7523) );
  OAI21X1 U18252 ( .A0(n3494), .A1(n7774), .B0(n7773), .Y(n7778) );
  OAI21X1 U18253 ( .A0(n7382), .A1(n26003), .B0(n6264), .Y(M0_a_8_) );
  XNOR2X1 U18254 ( .A(n15968), .B(n3196), .Y(n16126) );
  XNOR2X1 U18255 ( .A(n12519), .B(n12271), .Y(n12121) );
  XNOR2X1 U18256 ( .A(n12519), .B(n12561), .Y(n11688) );
  XNOR2X2 U18257 ( .A(n18902), .B(n18901), .Y(n23460) );
  XNOR2X1 U18258 ( .A(n17039), .B(n16884), .Y(n16127) );
  OAI22X1 U18259 ( .A0(n17060), .A1(n16201), .B0(n17061), .B1(n16241), .Y(
        n16251) );
  XNOR2X1 U18260 ( .A(n17039), .B(n3190), .Y(n16164) );
  OAI22X1 U18261 ( .A0(n6209), .A1(n15942), .B0(n25908), .B1(n25813), .Y(
        n11494) );
  ADDFHX4 U18262 ( .A(n12484), .B(n12483), .CI(n12482), .CO(n12494), .S(n12493) );
  NAND2X1 U18263 ( .A(n25229), .B(target_temp[22]), .Y(n11546) );
  OAI222X1 U18264 ( .A0(n26542), .A1(n23884), .B0(n3121), .B1(n24115), .C0(
        n4586), .C1(n24481), .Y(n2613) );
  OAI21XL U18265 ( .A0(n25731), .A1(n3121), .B0(n25730), .Y(n2574) );
  OAI22X1 U18266 ( .A0(n13576), .A1(n14157), .B0(n13619), .B1(n14120), .Y(
        n13632) );
  OAI22X1 U18267 ( .A0(n17148), .A1(n3190), .B0(n17147), .B1(n12561), .Y(
        n16936) );
  AOI22XL U18268 ( .A0(n24237), .A1(n23794), .B0(n2984), .B1(temp1[17]), .Y(
        n20675) );
  OAI21XL U18269 ( .A0(n10656), .A1(n10590), .B0(n10589), .Y(n10595) );
  OAI21XL U18270 ( .A0(n25813), .A1(n25913), .B0(n6190), .Y(n11484) );
  XNOR2X1 U18271 ( .A(n9886), .B(n9836), .Y(n9976) );
  XNOR2X1 U18272 ( .A(n3211), .B(n12561), .Y(n16124) );
  AND3X1 U18273 ( .A(n7885), .B(n26213), .C(n25886), .Y(n6174) );
  XNOR2X1 U18274 ( .A(n17264), .B(n17263), .Y(n6175) );
  AND2XL U18275 ( .A(n6568), .B(n6566), .Y(n6176) );
  XNOR2X1 U18276 ( .A(n18735), .B(n18734), .Y(n6182) );
  NAND2X4 U18277 ( .A(n13509), .B(n14291), .Y(n6191) );
  OAI21XL U18278 ( .A0(n26184), .A1(n21256), .B0(n21173), .Y(n21809) );
  OAI21XL U18279 ( .A0(n26177), .A1(n21256), .B0(n21235), .Y(n21862) );
  OAI21XL U18280 ( .A0(n26169), .A1(n21311), .B0(n21310), .Y(n21997) );
  OAI21XL U18281 ( .A0(n26173), .A1(n21256), .B0(n21247), .Y(n21901) );
  AND2XL U18282 ( .A(n16634), .B(n16633), .Y(n6197) );
  OAI21XL U18283 ( .A0(n26178), .A1(n21256), .B0(n21237), .Y(n21852) );
  OAI21XL U18284 ( .A0(n26179), .A1(n21331), .B0(n21240), .Y(n21844) );
  AND2XL U18285 ( .A(n9910), .B(n9909), .Y(n6201) );
  OAI21X2 U18286 ( .A0(n15558), .A1(n14875), .B0(n14920), .Y(n23966) );
  OAI21XL U18287 ( .A0(n26182), .A1(n21331), .B0(n21213), .Y(n21578) );
  OAI21XL U18288 ( .A0(n26175), .A1(n21256), .B0(n21254), .Y(n21875) );
  OAI21XL U18289 ( .A0(n26174), .A1(n21256), .B0(n21249), .Y(n21880) );
  OAI21XL U18290 ( .A0(n26176), .A1(n21256), .B0(n21252), .Y(n21870) );
  AND2XL U18291 ( .A(n13111), .B(n13110), .Y(n6204) );
  OR2XL U18292 ( .A(M2_b_19_), .B(M2_b_17_), .Y(n6206) );
  OAI21XL U18293 ( .A0(n26171), .A1(n21333), .B0(n21299), .Y(n21977) );
  AND2X2 U18294 ( .A(n6279), .B(n6231), .Y(n6469) );
  OR2X2 U18295 ( .A(n21759), .B(n21758), .Y(n6216) );
  OAI21X2 U18296 ( .A0(n21519), .A1(n21355), .B0(n21400), .Y(n23409) );
  AOI2BB1X2 U18297 ( .A0N(n22152), .A1N(n22258), .B0(n22213), .Y(n22188) );
  AND2X4 U18298 ( .A(n23967), .B(n26595), .Y(n6217) );
  INVX4 U18299 ( .A(n21429), .Y(n21519) );
  OAI21XL U18300 ( .A0(n26164), .A1(n21333), .B0(n21330), .Y(n21414) );
  OAI21XL U18301 ( .A0(n26163), .A1(n21333), .B0(n21316), .Y(n21410) );
  OAI21XL U18302 ( .A0(n26161), .A1(n21256), .B0(n21318), .Y(n21406) );
  OAI21XL U18303 ( .A0(n26165), .A1(n21333), .B0(n21323), .Y(n21435) );
  BUFX3 U18304 ( .A(n11493), .Y(M3_mult_x_15_b_12_) );
  AOI21XL U18305 ( .A0(n11140), .A1(n11395), .B0(n23089), .Y(n11142) );
  XOR2XL U18306 ( .A(n10768), .B(n11209), .Y(n10845) );
  XOR2XL U18307 ( .A(n10766), .B(n3054), .Y(n10867) );
  XOR2XL U18308 ( .A(n10801), .B(n3221), .Y(n10883) );
  XOR2XL U18309 ( .A(n23007), .B(n3055), .Y(n23017) );
  XOR2XL U18310 ( .A(n22968), .B(n3055), .Y(n23009) );
  XNOR2X1 U18311 ( .A(n3047), .B(n3110), .Y(n16629) );
  XOR2XL U18312 ( .A(n22608), .B(n3221), .Y(M6_mult_x_15_n1205) );
  XNOR2X1 U18313 ( .A(n16614), .B(n12271), .Y(n16594) );
  XNOR2XL U18314 ( .A(n25865), .B(n13204), .Y(n13113) );
  XOR2XL U18315 ( .A(n22690), .B(n3053), .Y(M6_mult_x_15_n1179) );
  XOR2XL U18316 ( .A(n22752), .B(n3054), .Y(M6_mult_x_15_n1153) );
  XNOR2XL U18317 ( .A(n18150), .B(n2978), .Y(n18152) );
  XNOR2X1 U18318 ( .A(n9904), .B(n9839), .Y(n9982) );
  AOI21XL U18319 ( .A0(n10900), .A1(n10899), .B0(n10898), .Y(n10903) );
  XOR2XL U18320 ( .A(n22744), .B(n3056), .Y(M6_mult_x_15_n1103) );
  OAI22XL U18321 ( .A0(n7093), .A1(n6406), .B0(n6365), .B1(n7094), .Y(n6404)
         );
  XNOR2XL U18322 ( .A(n4567), .B(n13204), .Y(n13157) );
  OAI22X1 U18323 ( .A0(n13209), .A1(n13972), .B0(n13172), .B1(n13971), .Y(
        n13213) );
  AOI21XL U18324 ( .A0(n22762), .A1(n22761), .B0(n22760), .Y(n22767) );
  XNOR2X1 U18325 ( .A(n9841), .B(n9863), .Y(n9753) );
  OAI22XL U18326 ( .A0(n9963), .A1(n9962), .B0(n9961), .B1(n3180), .Y(n9971)
         );
  XOR2XL U18327 ( .A(n22769), .B(n3054), .Y(M6_mult_x_15_n1150) );
  AOI21XL U18328 ( .A0(n6588), .A1(n6584), .B0(n6587), .Y(n6596) );
  XNOR2X1 U18329 ( .A(n12265), .B(n3190), .Y(n12117) );
  XNOR2XL U18330 ( .A(n18453), .B(n2978), .Y(n18042) );
  XNOR2X1 U18331 ( .A(n18503), .B(n2974), .Y(n18026) );
  XOR2XL U18332 ( .A(n22801), .B(n3221), .Y(M6_mult_x_15_n1197) );
  XOR2XL U18333 ( .A(n10853), .B(n10776), .Y(n22993) );
  XOR2XL U18334 ( .A(n10816), .B(n10815), .Y(n22998) );
  CLKINVX2 U18335 ( .A(n11166), .Y(n22989) );
  AOI22X1 U18336 ( .A0(n25229), .A1(y12[11]), .B0(n14427), .B1(y10[11]), .Y(
        n9202) );
  XNOR2XL U18337 ( .A(n23221), .B(n7621), .Y(n7197) );
  OAI21XL U18338 ( .A0(n3041), .A1(n19933), .B0(n19429), .Y(n19643) );
  OAI21XL U18339 ( .A0(n19929), .A1(n19747), .B0(n19547), .Y(n19548) );
  XOR2XL U18340 ( .A(n22738), .B(n3056), .Y(M6_mult_x_15_n1099) );
  XNOR2XL U18341 ( .A(n14357), .B(n14030), .Y(n13975) );
  XNOR2X1 U18342 ( .A(n10494), .B(n10342), .Y(n9464) );
  XOR2XL U18343 ( .A(n22850), .B(n3056), .Y(M6_mult_x_15_n1093) );
  XNOR2X1 U18344 ( .A(M2_mult_x_15_n43), .B(n9839), .Y(n9402) );
  AOI21XL U18345 ( .A0(n9933), .A1(n9929), .B0(n9932), .Y(n9942) );
  XNOR2X1 U18346 ( .A(n3199), .B(n16884), .Y(n16047) );
  OAI22X1 U18347 ( .A0(n7093), .A1(n3209), .B0(n7094), .B1(n26488), .Y(n7097)
         );
  OAI22X1 U18348 ( .A0(n7633), .A1(n7459), .B0(n7497), .B1(n7634), .Y(n7499)
         );
  XNOR2XL U18349 ( .A(n23219), .B(n25877), .Y(n7530) );
  XNOR2XL U18350 ( .A(n14266), .B(n25861), .Y(n13793) );
  OAI22X1 U18351 ( .A0(n13367), .A1(n14208), .B0(n13448), .B1(n14198), .Y(
        n13432) );
  XNOR2XL U18352 ( .A(n14028), .B(n14228), .Y(n13616) );
  XNOR2X1 U18353 ( .A(n25864), .B(n4848), .Y(n13601) );
  XNOR2X1 U18354 ( .A(M3_mult_x_15_a_17_), .B(n12271), .Y(n12005) );
  XNOR2X1 U18355 ( .A(n18500), .B(n3049), .Y(n17942) );
  AOI21XL U18356 ( .A0(n21638), .A1(n3222), .B0(n21849), .Y(n21637) );
  AOI21XL U18357 ( .A0(n21851), .A1(n3222), .B0(n21849), .Y(n21850) );
  NOR2X1 U18358 ( .A(n14875), .B(n14946), .Y(n14878) );
  XOR2XL U18359 ( .A(n22750), .B(n3056), .Y(M6_mult_x_15_n1088) );
  XOR2XL U18360 ( .A(n21075), .B(n3058), .Y(M6_mult_x_15_n1058) );
  XOR2XL U18361 ( .A(n22735), .B(n3054), .Y(M6_mult_x_15_n1141) );
  XOR2XL U18362 ( .A(n22624), .B(n3221), .Y(M6_mult_x_15_n1195) );
  XOR2XL U18363 ( .A(n22790), .B(n3054), .Y(M6_mult_x_15_n1143) );
  XOR2XL U18364 ( .A(n22900), .B(n3221), .Y(M6_mult_x_15_n1193) );
  OAI22X1 U18365 ( .A0(n13840), .A1(n13972), .B0(n13777), .B1(n13971), .Y(
        n13846) );
  XNOR2XL U18366 ( .A(n14195), .B(n23173), .Y(n14071) );
  XNOR2XL U18367 ( .A(n14235), .B(M1_b_19_), .Y(n14069) );
  OAI22X1 U18368 ( .A0(n10660), .A1(n9863), .B0(n3178), .B1(n9836), .Y(n9466)
         );
  OAI22X1 U18369 ( .A0(n2993), .A1(n14117), .B0(n14289), .B1(n14196), .Y(
        n14091) );
  OAI22X1 U18370 ( .A0(n9504), .A1(n9340), .B0(n10496), .B1(n9460), .Y(n9470)
         );
  OAI22XL U18371 ( .A0(n9551), .A1(n9295), .B0(n9838), .B1(n9227), .Y(n9263)
         );
  XNOR2X1 U18372 ( .A(n3022), .B(n3190), .Y(n16318) );
  NOR2X1 U18373 ( .A(n19901), .B(n19437), .Y(n19245) );
  AOI21XL U18374 ( .A0(n15125), .A1(n23955), .B0(n15573), .Y(n15124) );
  XNOR2X1 U18375 ( .A(n12594), .B(n3190), .Y(n11811) );
  XNOR2X1 U18376 ( .A(n12716), .B(n3197), .Y(n11722) );
  OAI21XL U18377 ( .A0(n19566), .A1(n19923), .B0(n19446), .Y(n19625) );
  OAI21XL U18378 ( .A0(n3165), .A1(n19507), .B0(n19506), .Y(n19767) );
  OAI21XL U18379 ( .A0(n26168), .A1(n21311), .B0(n21292), .Y(n21987) );
  AOI21XL U18380 ( .A0(n8685), .A1(n8823), .B0(n3155), .Y(n8684) );
  XOR2XL U18381 ( .A(n22503), .B(n3058), .Y(M6_mult_x_15_n1062) );
  XOR2XL U18382 ( .A(n21061), .B(n3058), .Y(M6_mult_x_15_n1056) );
  OAI22X1 U18383 ( .A0(n12759), .A1(n11690), .B0(n12760), .B1(n11689), .Y(
        n11701) );
  OAI22X1 U18384 ( .A0(n12597), .A1(n11842), .B0(n12595), .B1(n11811), .Y(
        n11857) );
  XNOR2XL U18385 ( .A(n12716), .B(M3_mult_x_15_b_19_), .Y(n12516) );
  XNOR2XL U18386 ( .A(n18804), .B(n18803), .Y(n18805) );
  OAI22X1 U18387 ( .A0(n18624), .A1(n17507), .B0(n18625), .B1(n17506), .Y(
        n17566) );
  OAI21XL U18388 ( .A0(n8645), .A1(n8926), .B0(n8644), .Y(n8917) );
  AOI21XL U18389 ( .A0(n8538), .A1(n8592), .B0(n8536), .Y(n8541) );
  OAI21XL U18390 ( .A0(n15392), .A1(n15676), .B0(n15391), .Y(n15667) );
  AOI21XL U18391 ( .A0(n7952), .A1(n7951), .B0(n7950), .Y(n7953) );
  NOR2X1 U18392 ( .A(n18941), .B(n18951), .Y(n18690) );
  AOI21XL U18393 ( .A0(n14534), .A1(n14539), .B0(n14485), .Y(n14486) );
  AOI21XL U18394 ( .A0(n22020), .A1(n22060), .B0(n22019), .Y(n22021) );
  XOR2XL U18395 ( .A(n11123), .B(n11122), .Y(n11462) );
  AOI21XL U18396 ( .A0(n11390), .A1(n11389), .B0(n11388), .Y(n11391) );
  AOI21XL U18397 ( .A0(n19961), .A1(n20001), .B0(n19960), .Y(n19962) );
  AOI21XL U18398 ( .A0(n15582), .A1(n15622), .B0(n15581), .Y(n15583) );
  XOR2X1 U18399 ( .A(n22092), .B(n22091), .Y(n22305) );
  XOR2XL U18400 ( .A(n11045), .B(n11027), .Y(n20625) );
  AOI21XL U18401 ( .A0(n3072), .A1(n24893), .B0(n24892), .Y(n24897) );
  XOR2XL U18402 ( .A(n23500), .B(n23499), .Y(n23946) );
  XOR2XL U18403 ( .A(n23470), .B(n23469), .Y(n23726) );
  OAI21XL U18404 ( .A0(n19564), .A1(n19321), .B0(n19320), .Y(n23204) );
  AOI21XL U18405 ( .A0(n25013), .A1(n25012), .B0(n15688), .Y(n25014) );
  OAI21XL U18406 ( .A0(n21519), .A1(n21416), .B0(n21415), .Y(n23119) );
  XOR2XL U18407 ( .A(n20295), .B(n20294), .Y(n20627) );
  XOR2XL U18408 ( .A(n20768), .B(n20767), .Y(n20824) );
  XOR2XL U18409 ( .A(n9174), .B(n9173), .Y(n20800) );
  XOR2XL U18410 ( .A(n11596), .B(n13013), .Y(n11612) );
  XOR2XL U18411 ( .A(n14449), .B(n14701), .Y(n14464) );
  AOI21XL U18412 ( .A0(n22406), .A1(n3079), .B0(n22405), .Y(n23270) );
  AOI21XL U18413 ( .A0(n24012), .A1(n24013), .B0(n23984), .Y(n23986) );
  XOR2XL U18414 ( .A(n23684), .B(n23685), .Y(n23686) );
  XOR2XL U18415 ( .A(n17180), .B(n17402), .Y(n17194) );
  XOR2XL U18416 ( .A(n21168), .B(n22484), .Y(n21169) );
  OAI21XL U18417 ( .A0(n25531), .A1(n3121), .B0(n23931), .Y(n2600) );
  OAI21XL U18418 ( .A0(n25747), .A1(n3121), .B0(n20732), .Y(n2572) );
  OAI21XL U18419 ( .A0(mul5_out[23]), .A1(n5434), .B0(n25223), .Y(n2342) );
  OAI21XL U18420 ( .A0(n25577), .A1(n25584), .B0(n25576), .Y(n2025) );
  OAI21XL U18421 ( .A0(n25712), .A1(n25711), .B0(n25710), .Y(n2160) );
  OAI21XL U18422 ( .A0(n25508), .A1(n4572), .B0(n25507), .Y(n2049) );
  CLKINVX4 U18423 ( .A(n6476), .Y(n25868) );
  AOI21X1 U18424 ( .A0(n6733), .A1(y10[10]), .B0(n25148), .Y(n6226) );
  NOR2X1 U18425 ( .A(n4583), .B(n6227), .Y(n25147) );
  OAI21XL U18426 ( .A0(n6274), .A1(n26214), .B0(n6228), .Y(M0_b_10_) );
  INVX1 U18427 ( .A(M0_a_0_), .Y(n6231) );
  BUFX3 U18428 ( .A(M0_b_18_), .Y(n25875) );
  AOI22XL U18429 ( .A0(n7389), .A1(target_temp[19]), .B0(in_valid_d), .B1(
        w1[19]), .Y(n6232) );
  AOI21XL U18430 ( .A0(n6733), .A1(y10[2]), .B0(n25140), .Y(n6234) );
  INVX4 U18431 ( .A(n7644), .Y(n25870) );
  AOI22XL U18432 ( .A0(n7389), .A1(target_temp[8]), .B0(in_valid_d), .B1(w1[8]), .Y(n6240) );
  OAI21XL U18433 ( .A0(n6274), .A1(n26220), .B0(n6240), .Y(M0_b_8_) );
  OAI21XL U18434 ( .A0(n6274), .A1(n26226), .B0(n6241), .Y(M0_b_0_) );
  NOR2X1 U18435 ( .A(n4586), .B(n6242), .Y(n25143) );
  AOI21XL U18436 ( .A0(n6733), .A1(y10[6]), .B0(n25144), .Y(n6245) );
  AOI22XL U18437 ( .A0(n7389), .A1(target_temp[11]), .B0(in_valid_d), .B1(
        w1[11]), .Y(n6248) );
  AOI22XL U18438 ( .A0(n7389), .A1(target_temp[5]), .B0(in_valid_d), .B1(w1[5]), .Y(n6251) );
  AOI22XL U18439 ( .A0(n7389), .A1(target_temp[15]), .B0(in_valid_d), .B1(
        w1[15]), .Y(n6253) );
  AOI22XL U18440 ( .A0(n7389), .A1(target_temp[7]), .B0(in_valid_d), .B1(w1[7]), .Y(n6254) );
  OAI21XL U18441 ( .A0(n6274), .A1(n26219), .B0(n6254), .Y(M0_b_7_) );
  OAI21X1 U18442 ( .A0(n7382), .A1(n26016), .B0(n6256), .Y(M0_a_20_) );
  OAI21XL U18443 ( .A0(n6274), .A1(n26230), .B0(n6257), .Y(M0_b_20_) );
  CLKINVX3 U18444 ( .A(M0_a_15_), .Y(n7564) );
  BUFX3 U18445 ( .A(M0_b_15_), .Y(n25877) );
  NOR2X1 U18446 ( .A(n4583), .B(n6263), .Y(n25146) );
  AOI21XL U18447 ( .A0(n6733), .A1(y10[8]), .B0(n25146), .Y(n6264) );
  AOI21XL U18448 ( .A0(n6733), .A1(y10[16]), .B0(n25154), .Y(n6268) );
  AOI22XL U18449 ( .A0(n6733), .A1(target_temp[21]), .B0(in_valid_d), .B1(
        w1[21]), .Y(n6272) );
  AOI22XL U18450 ( .A0(n6733), .A1(target_temp[22]), .B0(in_valid_d), .B1(
        w1[22]), .Y(n6273) );
  NAND2X4 U18451 ( .A(n23970), .B(cs[2]), .Y(n26595) );
  XNOR2XL U18452 ( .A(M0_b_9_), .B(n25868), .Y(n6283) );
  XOR2X1 U18453 ( .A(n7220), .B(M0_a_10_), .Y(n6276) );
  INVX8 U18454 ( .A(n6275), .Y(n7512) );
  NAND2X4 U18455 ( .A(n6276), .B(n7512), .Y(n7511) );
  XNOR2X1 U18456 ( .A(n25868), .B(n25880), .Y(n6758) );
  OAI22XL U18457 ( .A0(n6283), .A1(n7511), .B0(n7512), .B1(n6758), .Y(n6761)
         );
  NOR2X1 U18458 ( .A(n4586), .B(n6277), .Y(n25139) );
  OAI21X1 U18459 ( .A0(n7382), .A1(n25997), .B0(n6278), .Y(n6279) );
  INVX4 U18460 ( .A(n6469), .Y(n6845) );
  CLKINVX3 U18461 ( .A(n6279), .Y(n6861) );
  CLKINVX3 U18462 ( .A(n6861), .Y(n6928) );
  CLKINVX4 U18463 ( .A(n6861), .Y(n21054) );
  OAI22XL U18464 ( .A0(n6845), .A1(n6284), .B0(n6290), .B1(n6843), .Y(n6344)
         );
  XNOR2XL U18465 ( .A(n25866), .B(n6830), .Y(n6286) );
  XNOR2XL U18466 ( .A(M0_b_1_), .B(n25870), .Y(n6346) );
  AOI21XL U18467 ( .A0(n6733), .A1(y10[17]), .B0(n25155), .Y(n6280) );
  XOR2X4 U18468 ( .A(n6299), .B(n6281), .Y(n7695) );
  XNOR2XL U18469 ( .A(M0_b_2_), .B(n25870), .Y(n6784) );
  XNOR2X1 U18470 ( .A(n25868), .B(n7475), .Y(n6287) );
  INVXL U18471 ( .A(M0_b_0_), .Y(n6324) );
  XNOR2X1 U18472 ( .A(n21054), .B(n7646), .Y(n6321) );
  OAI22X1 U18473 ( .A0(n6845), .A1(n6321), .B0(n6284), .B1(n6231), .Y(n6332)
         );
  XNOR2X1 U18474 ( .A(n25867), .B(n25879), .Y(n6322) );
  XNOR2X1 U18475 ( .A(n25867), .B(n7569), .Y(n6296) );
  OAI22XL U18476 ( .A0(n6613), .A1(n6322), .B0(n7146), .B1(n6296), .Y(n6331)
         );
  XNOR2X1 U18477 ( .A(n23220), .B(n7164), .Y(n6301) );
  XNOR2X1 U18478 ( .A(n23220), .B(n25882), .Y(n6312) );
  XNOR2XL U18479 ( .A(n25866), .B(M0_b_15_), .Y(n6302) );
  OAI22XL U18480 ( .A0(n7511), .A1(n6303), .B0(n7512), .B1(n6287), .Y(n6305)
         );
  XNOR2X1 U18481 ( .A(n6288), .B(M0_a_20_), .Y(n6289) );
  NOR2BX1 U18482 ( .AN(n6944), .B(n7712), .Y(n6787) );
  XNOR2X1 U18483 ( .A(n21054), .B(n25873), .Y(n6749) );
  OAI22X1 U18484 ( .A0(n6845), .A1(n6290), .B0(n6749), .B1(n6843), .Y(n6786)
         );
  XNOR2X1 U18485 ( .A(n25869), .B(n7164), .Y(n6313) );
  XNOR2XL U18486 ( .A(n25869), .B(M0_b_6_), .Y(n6737) );
  OAI22XL U18487 ( .A0(n4592), .A1(n6313), .B0(n3046), .B1(n6737), .Y(n6785)
         );
  XNOR2X1 U18488 ( .A(n3209), .B(n25877), .Y(n6340) );
  INVX4 U18489 ( .A(n6293), .Y(n7094) );
  XNOR2XL U18490 ( .A(n7286), .B(n25880), .Y(n6304) );
  XNOR2X1 U18491 ( .A(n7286), .B(n25879), .Y(n6297) );
  INVX4 U18492 ( .A(n6295), .Y(n7288) );
  OAI22X1 U18493 ( .A0(n7287), .A1(n6304), .B0(n6297), .B1(n7288), .Y(n6309)
         );
  XNOR2X1 U18494 ( .A(n25867), .B(n25878), .Y(n6342) );
  OAI22XL U18495 ( .A0(n6613), .A1(n6296), .B0(n6608), .B1(n6342), .Y(n6308)
         );
  XNOR2XL U18496 ( .A(n7286), .B(n7569), .Y(n6756) );
  OAI22XL U18497 ( .A0(n7287), .A1(n6297), .B0(n6756), .B1(n7288), .Y(n6755)
         );
  XNOR2X1 U18498 ( .A(n23220), .B(n25881), .Y(n6311) );
  XNOR2X1 U18499 ( .A(n23220), .B(n7475), .Y(n6751) );
  XNOR2X1 U18500 ( .A(n23221), .B(n7165), .Y(n6757) );
  OAI22XL U18501 ( .A0(n6348), .A1(n7633), .B0(n6757), .B1(n7634), .Y(n6753)
         );
  XNOR2X1 U18502 ( .A(n23220), .B(n7165), .Y(n6377) );
  OAI22XL U18503 ( .A0(n7535), .A1(n6377), .B0(n6301), .B1(n7460), .Y(n6370)
         );
  XNOR2XL U18504 ( .A(n25866), .B(n7621), .Y(n6367) );
  OAI22XL U18505 ( .A0(n7511), .A1(n6363), .B0(n7512), .B1(n6303), .Y(n6368)
         );
  XNOR2X1 U18506 ( .A(n25869), .B(n7165), .Y(n6314) );
  XNOR2X1 U18507 ( .A(n3209), .B(n25878), .Y(n6319) );
  XNOR2XL U18508 ( .A(M0_b_9_), .B(n4789), .Y(n6323) );
  OAI22XL U18509 ( .A0(n6323), .A1(n7287), .B0(n6304), .B1(n7288), .Y(n6316)
         );
  CMPR32X1 U18510 ( .A(n6307), .B(n6306), .C(n6305), .CO(n6356), .S(n6371) );
  OAI22XL U18511 ( .A0(n7093), .A1(n6365), .B0(n6319), .B1(n7094), .Y(n6376)
         );
  XNOR2X1 U18512 ( .A(n25867), .B(n25880), .Y(n6393) );
  XNOR2XL U18513 ( .A(n7286), .B(M0_b_8_), .Y(n6364) );
  XNOR2XL U18514 ( .A(n23221), .B(n6944), .Y(n6325) );
  XNOR2X1 U18515 ( .A(M0_b_2_), .B(n25869), .Y(n6380) );
  OAI22XL U18516 ( .A0(n6380), .A1(n4592), .B0(n6327), .B1(n3046), .Y(n6381)
         );
  ADDHXL U18517 ( .A(n6329), .B(n6328), .CO(n6355), .S(n6374) );
  XNOR2XL U18518 ( .A(M0_b_2_), .B(n23221), .Y(n6349) );
  XNOR2X1 U18519 ( .A(n3209), .B(n25876), .Y(n6734) );
  OAI22XL U18520 ( .A0(n7093), .A1(n6340), .B0(n6734), .B1(n7094), .Y(n6740)
         );
  XNOR2X1 U18521 ( .A(n25866), .B(n25875), .Y(n6750) );
  OAI22X1 U18522 ( .A0(n6991), .A1(n6341), .B0(n6990), .B1(n6750), .Y(n6739)
         );
  OAI22XL U18523 ( .A0(n6613), .A1(n6342), .B0(n6608), .B1(n6735), .Y(n6738)
         );
  OAI22XL U18524 ( .A0(n6349), .A1(n7633), .B0(n6348), .B1(n6300), .Y(n6350)
         );
  ADDFHX1 U18525 ( .A(n6352), .B(n6351), .CI(n6350), .CO(n6798), .S(n6361) );
  ADDFHX1 U18526 ( .A(n6355), .B(n6354), .CI(n6353), .CO(n6360), .S(n6390) );
  ADDFHX1 U18527 ( .A(n6361), .B(n6360), .CI(n6359), .CO(n6804), .S(n6389) );
  XNOR2X1 U18528 ( .A(n21054), .B(n25877), .Y(n6378) );
  OAI22X1 U18529 ( .A0(n6845), .A1(n6378), .B0(n6362), .B1(n6843), .Y(n6395)
         );
  XNOR2X1 U18530 ( .A(n25868), .B(n7164), .Y(n6379) );
  OAI22XL U18531 ( .A0(n7511), .A1(n6379), .B0(n7512), .B1(n6363), .Y(n6394)
         );
  XNOR2X1 U18532 ( .A(n4789), .B(n25881), .Y(n6397) );
  XNOR2X1 U18533 ( .A(n3209), .B(n25879), .Y(n6406) );
  XNOR2XL U18534 ( .A(n25866), .B(n25878), .Y(n6399) );
  OAI22XL U18535 ( .A0(n6991), .A1(n6399), .B0(n6602), .B1(n6367), .Y(n6403)
         );
  ADDFHX1 U18536 ( .A(n6370), .B(n6369), .CI(n6368), .CO(n6373), .S(n6400) );
  CMPR32X1 U18537 ( .A(n6376), .B(n6375), .C(n6374), .CO(n6392), .S(n6423) );
  OAI22XL U18538 ( .A0(n6425), .A1(n7535), .B0(n6377), .B1(n7460), .Y(n6413)
         );
  XNOR2X1 U18539 ( .A(n21054), .B(n7621), .Y(n6426) );
  OAI22XL U18540 ( .A0(n6845), .A1(n6426), .B0(n6378), .B1(n6843), .Y(n6408)
         );
  XNOR2X1 U18541 ( .A(n25868), .B(n7165), .Y(n6433) );
  OAI22XL U18542 ( .A0(n6410), .A1(n4592), .B0(n6380), .B1(n3046), .Y(n6411)
         );
  XNOR2X1 U18543 ( .A(M0_b_9_), .B(n25867), .Y(n6424) );
  OAI22XL U18544 ( .A0(n6424), .A1(n6613), .B0(n6608), .B1(n6393), .Y(n6430)
         );
  ADDFHX1 U18545 ( .A(n6396), .B(n6395), .CI(n6394), .CO(n6402), .S(n6429) );
  OAI22XL U18546 ( .A0(n7287), .A1(n6431), .B0(n6397), .B1(n7288), .Y(n6436)
         );
  XNOR2XL U18547 ( .A(n25866), .B(n7569), .Y(n6427) );
  OAI22XL U18548 ( .A0(n6991), .A1(n6427), .B0(n6602), .B1(n6399), .Y(n6434)
         );
  OAI22XL U18549 ( .A0(n7093), .A1(n6449), .B0(n6406), .B1(n7094), .Y(n6439)
         );
  CMPR22X1 U18550 ( .A(n4736), .B(n6407), .CO(n6412), .S(n6438) );
  OAI22XL U18551 ( .A0(n6410), .A1(n3046), .B0(n4592), .B1(n6409), .Y(n6437)
         );
  ADDFHX1 U18552 ( .A(n6413), .B(n6412), .CI(n6411), .CO(n6422), .S(n6446) );
  ADDFHX1 U18553 ( .A(n6420), .B(n6418), .CI(n6419), .CO(n6729), .S(n6726) );
  ADDFHX1 U18554 ( .A(n6423), .B(n6422), .CI(n6421), .CO(n6414), .S(n6445) );
  XNOR2X1 U18555 ( .A(n25867), .B(n7475), .Y(n6432) );
  OAI22XL U18556 ( .A0(n6424), .A1(n6608), .B0(n6613), .B1(n6432), .Y(n6455)
         );
  XNOR2XL U18557 ( .A(M0_b_2_), .B(n23220), .Y(n6452) );
  OAI22XL U18558 ( .A0(n6452), .A1(n7535), .B0(n6425), .B1(n7460), .Y(n6454)
         );
  XNOR2X1 U18559 ( .A(n21054), .B(n25878), .Y(n6450) );
  OAI22XL U18560 ( .A0(n6845), .A1(n6450), .B0(n6426), .B1(n6231), .Y(n6457)
         );
  XNOR2XL U18561 ( .A(n25866), .B(n25879), .Y(n6461) );
  OAI22XL U18562 ( .A0(n6991), .A1(n6461), .B0(n6602), .B1(n6427), .Y(n6456)
         );
  XNOR2X1 U18563 ( .A(n4789), .B(n7164), .Y(n6459) );
  OAI22XL U18564 ( .A0(n7287), .A1(n6459), .B0(n6431), .B1(n7288), .Y(n6464)
         );
  XNOR2X1 U18565 ( .A(n25867), .B(n25881), .Y(n6451) );
  OAI22X1 U18566 ( .A0(n6613), .A1(n6451), .B0(n6608), .B1(n6432), .Y(n6463)
         );
  XNOR2XL U18567 ( .A(n4806), .B(n25868), .Y(n6541) );
  OAI22XL U18568 ( .A0(n6541), .A1(n7511), .B0(n7512), .B1(n6433), .Y(n6462)
         );
  ADDFHX1 U18569 ( .A(n6439), .B(n6438), .CI(n6437), .CO(n6447), .S(n6694) );
  ADDFHX1 U18570 ( .A(n6442), .B(n6441), .CI(n6440), .CO(n6419), .S(n6443) );
  ADDFHX1 U18571 ( .A(n6445), .B(n6444), .CI(n6443), .CO(n6725), .S(n6723) );
  XNOR2X1 U18572 ( .A(M0_b_9_), .B(n3209), .Y(n6524) );
  OAI22XL U18573 ( .A0(n6524), .A1(n7093), .B0(n6449), .B1(n7094), .Y(n6687)
         );
  XNOR2X1 U18574 ( .A(n21054), .B(n7569), .Y(n6470) );
  XNOR2X1 U18575 ( .A(n25867), .B(n25882), .Y(n6472) );
  OAI22X1 U18576 ( .A0(n6613), .A1(n6472), .B0(n6608), .B1(n6451), .Y(n6537)
         );
  XNOR2XL U18577 ( .A(M0_b_1_), .B(n23220), .Y(n6540) );
  OAI22XL U18578 ( .A0(n6540), .A1(n7535), .B0(n6452), .B1(n7460), .Y(n6685)
         );
  XNOR2X1 U18579 ( .A(n4789), .B(n7165), .Y(n6486) );
  OAI22XL U18580 ( .A0(n7287), .A1(n6486), .B0(n6459), .B1(n7288), .Y(n6530)
         );
  OAI22XL U18581 ( .A0(n7535), .A1(n7534), .B0(n7460), .B1(n6460), .Y(n6529)
         );
  XNOR2XL U18582 ( .A(n25866), .B(M0_b_10_), .Y(n6485) );
  OAI22XL U18583 ( .A0(n6991), .A1(n6485), .B0(n6602), .B1(n6461), .Y(n6528)
         );
  XNOR2X1 U18584 ( .A(n21054), .B(n25880), .Y(n6497) );
  OAI22XL U18585 ( .A0(n6845), .A1(n6497), .B0(n6471), .B1(n6843), .Y(n6478)
         );
  XNOR2X1 U18586 ( .A(n25867), .B(n7164), .Y(n6473) );
  OAI22XL U18587 ( .A0(n6613), .A1(n6479), .B0(n6608), .B1(n6473), .Y(n6477)
         );
  XNOR2XL U18588 ( .A(M0_b_1_), .B(n25868), .Y(n6489) );
  XNOR2XL U18589 ( .A(M0_b_2_), .B(n25868), .Y(n6542) );
  OAI22XL U18590 ( .A0(n6613), .A1(n6473), .B0(n6608), .B1(n6472), .Y(n6525)
         );
  XNOR2X1 U18591 ( .A(n7092), .B(n7164), .Y(n6500) );
  XNOR2XL U18592 ( .A(n25866), .B(n7475), .Y(n6490) );
  OAI22XL U18593 ( .A0(n7093), .A1(n6474), .B0(n6487), .B1(n7094), .Y(n6484)
         );
  ADDHXL U18594 ( .A(n6478), .B(n6477), .CO(n6545), .S(n6482) );
  OAI22XL U18595 ( .A0(n6515), .A1(n6613), .B0(n6608), .B1(n6479), .Y(n6512)
         );
  XNOR2XL U18596 ( .A(M0_b_1_), .B(n4789), .Y(n6503) );
  XNOR2XL U18597 ( .A(M0_b_2_), .B(n4789), .Y(n6493) );
  OAI22XL U18598 ( .A0(n7287), .A1(n3213), .B0(n7288), .B1(n6480), .Y(n6514)
         );
  XNOR2XL U18599 ( .A(n25866), .B(n25882), .Y(n6517) );
  OAI22XL U18600 ( .A0(n6991), .A1(n6517), .B0(n6602), .B1(n6481), .Y(n6513)
         );
  OAI22XL U18601 ( .A0(n6491), .A1(n6991), .B0(n6602), .B1(n6485), .Y(n6536)
         );
  XNOR2XL U18602 ( .A(n4806), .B(n4789), .Y(n6492) );
  OAI22XL U18603 ( .A0(n6492), .A1(n7287), .B0(n6486), .B1(n7288), .Y(n6535)
         );
  XNOR2XL U18604 ( .A(n3209), .B(n7475), .Y(n6523) );
  OAI22XL U18605 ( .A0(n7093), .A1(n6487), .B0(n6523), .B1(n7094), .Y(n6534)
         );
  XNOR2XL U18606 ( .A(n25868), .B(n6944), .Y(n6488) );
  OAI22XL U18607 ( .A0(n6489), .A1(n7512), .B0(n7511), .B1(n6488), .Y(n6496)
         );
  OAI22XL U18608 ( .A0(n6491), .A1(n6990), .B0(n6991), .B1(n6490), .Y(n6495)
         );
  OAI22XL U18609 ( .A0(n6493), .A1(n7287), .B0(n6492), .B1(n7288), .Y(n6494)
         );
  CMPR32X1 U18610 ( .A(n6496), .B(n6495), .C(n6494), .CO(n6531), .S(n6509) );
  XNOR2X1 U18611 ( .A(n7092), .B(n7165), .Y(n6609) );
  OAI22XL U18612 ( .A0(n7093), .A1(n6609), .B0(n6500), .B1(n7094), .Y(n6645)
         );
  XNOR2XL U18613 ( .A(n4789), .B(n6944), .Y(n6502) );
  OAI22XL U18614 ( .A0(n6503), .A1(n7288), .B0(n7287), .B1(n6502), .Y(n6643)
         );
  ADDFHX1 U18615 ( .A(n6506), .B(n6505), .CI(n6504), .CO(n6547), .S(n6507) );
  ADDHXL U18616 ( .A(n6514), .B(n6513), .CO(n6510), .S(n6651) );
  OAI22XL U18617 ( .A0(n6612), .A1(n6613), .B0(n6515), .B1(n7146), .Y(n6650)
         );
  XNOR2XL U18618 ( .A(n21054), .B(M0_b_7_), .Y(n6604) );
  OAI22XL U18619 ( .A0(n6845), .A1(n6604), .B0(n6516), .B1(n6843), .Y(n6599)
         );
  OAI22XL U18620 ( .A0(n6991), .A1(n6601), .B0(n6602), .B1(n6517), .Y(n6598)
         );
  NOR2XL U18621 ( .A(n6667), .B(n6666), .Y(n6521) );
  INVXL U18622 ( .A(n6521), .Y(n6522) );
  CMPR22X1 U18623 ( .A(n6538), .B(n6537), .CO(n6686), .S(n6684) );
  OAI22XL U18624 ( .A0(n6542), .A1(n7511), .B0(n6541), .B1(n7512), .Y(n6682)
         );
  ADDFHX1 U18625 ( .A(n6545), .B(n6544), .CI(n6543), .CO(n6679), .S(n6548) );
  ADDFHX1 U18626 ( .A(n6548), .B(n6547), .CI(n6546), .CO(n6672), .S(n6669) );
  XNOR2X1 U18627 ( .A(n21054), .B(n7165), .Y(n6560) );
  XNOR2X1 U18628 ( .A(n21054), .B(n7164), .Y(n6550) );
  OAI22XL U18629 ( .A0(n6845), .A1(n6560), .B0(n6550), .B1(n6843), .Y(n6552)
         );
  OAI22XL U18630 ( .A0(n7093), .A1(n26488), .B0(n7094), .B1(n6549), .Y(n6551)
         );
  OAI22XL U18631 ( .A0(n6845), .A1(n6550), .B0(n6605), .B1(n6843), .Y(n6618)
         );
  OAI22XL U18632 ( .A0(n6555), .A1(n6991), .B0(n6602), .B1(n6603), .Y(n6617)
         );
  ADDHXL U18633 ( .A(n6552), .B(n6551), .CO(n6628), .S(n6559) );
  XNOR2XL U18634 ( .A(n7092), .B(n6944), .Y(n6553) );
  XNOR2X1 U18635 ( .A(M0_b_2_), .B(n25866), .Y(n6561) );
  OAI22XL U18636 ( .A0(n6561), .A1(n6991), .B0(n6555), .B1(n6602), .Y(n6557)
         );
  ADDFHX1 U18637 ( .A(n6559), .B(n6558), .CI(n6557), .CO(n6591), .S(n6590) );
  NAND2XL U18638 ( .A(n6556), .B(n6562), .Y(n6597) );
  XNOR2XL U18639 ( .A(M0_b_2_), .B(n21054), .Y(n6573) );
  INVXL U18640 ( .A(n6563), .Y(n6564) );
  AND2XL U18641 ( .A(n6565), .B(n6564), .Y(n6567) );
  AOI21XL U18642 ( .A0(n6568), .A1(n6567), .B0(n6176), .Y(n6578) );
  OAI22X1 U18643 ( .A0(n6991), .A1(n6989), .B0(n6602), .B1(n6569), .Y(n6583)
         );
  XNOR2XL U18644 ( .A(n25866), .B(n6944), .Y(n6570) );
  OAI22X1 U18645 ( .A0(n6571), .A1(n6990), .B0(n6991), .B1(n6570), .Y(n6582)
         );
  NOR2XL U18646 ( .A(n6575), .B(n6574), .Y(n6577) );
  NAND2XL U18647 ( .A(n6575), .B(n6574), .Y(n6576) );
  OAI21XL U18648 ( .A0(n6578), .A1(n6577), .B0(n6576), .Y(n6588) );
  CMPR32X1 U18649 ( .A(n6581), .B(n6580), .C(n6579), .CO(n6589), .S(n6586) );
  CMPR22X1 U18650 ( .A(n6583), .B(n6582), .CO(n6585), .S(n6575) );
  AND2XL U18651 ( .A(n6586), .B(n6585), .Y(n6587) );
  AOI21XL U18652 ( .A0(n6556), .A1(n6594), .B0(n6593), .Y(n6595) );
  OAI21XL U18653 ( .A0(n6597), .A1(n6596), .B0(n6595), .Y(n6639) );
  OAI22XL U18654 ( .A0(n6991), .A1(n6603), .B0(n6602), .B1(n6601), .Y(n6622)
         );
  OAI22XL U18655 ( .A0(n6614), .A1(n6608), .B0(n6613), .B1(n6607), .Y(n6620)
         );
  OAI22XL U18656 ( .A0(n6615), .A1(n7093), .B0(n6609), .B1(n7094), .Y(n6648)
         );
  CMPR22X1 U18657 ( .A(n4738), .B(n6610), .CO(n6647), .S(n6621) );
  ADDFHX1 U18658 ( .A(n6622), .B(n6621), .CI(n6620), .CO(n6656), .S(n6623) );
  NOR2X1 U18659 ( .A(n6633), .B(n6632), .Y(n6636) );
  CMPR32X1 U18660 ( .A(n6625), .B(n6624), .C(n6623), .CO(n6632), .S(n6631) );
  NOR2XL U18661 ( .A(n6631), .B(n6630), .Y(n6629) );
  NOR2X1 U18662 ( .A(n6636), .B(n6629), .Y(n6638) );
  NAND2XL U18663 ( .A(n6631), .B(n6630), .Y(n6635) );
  NAND2XL U18664 ( .A(n6633), .B(n6632), .Y(n6634) );
  OAI21XL U18665 ( .A0(n6636), .A1(n6635), .B0(n6634), .Y(n6637) );
  AOI21XL U18666 ( .A0(n6639), .A1(n6638), .B0(n6637), .Y(n6665) );
  CMPR32X1 U18667 ( .A(n6642), .B(n6641), .C(n6640), .CO(n6666), .S(n6662) );
  ADDFHX1 U18668 ( .A(n6651), .B(n4760), .CI(n6649), .CO(n6641), .S(n6652) );
  CMPR32X1 U18669 ( .A(n6657), .B(n6656), .C(n6655), .CO(n6659), .S(n6633) );
  OR2X2 U18670 ( .A(n6660), .B(n6659), .Y(n6658) );
  NAND2XL U18671 ( .A(n6673), .B(n6672), .Y(n6674) );
  ADDFHX1 U18672 ( .A(n6678), .B(n6677), .CI(n6676), .CO(n6700), .S(n6705) );
  ADDFHX1 U18673 ( .A(n6681), .B(n6680), .CI(n6679), .CO(n6704), .S(n6691) );
  CMPR32X1 U18674 ( .A(n6705), .B(n6704), .C(n6703), .CO(n6714), .S(n6713) );
  ADDFHX1 U18675 ( .A(n6711), .B(n6710), .CI(n6709), .CO(n6718), .S(n6715) );
  XNOR2XL U18676 ( .A(M0_b_9_), .B(n23220), .Y(n6752) );
  XNOR2X1 U18677 ( .A(n23220), .B(n25880), .Y(n6819) );
  OAI22XL U18678 ( .A0(n6752), .A1(n7535), .B0(n6819), .B1(n7460), .Y(n6854)
         );
  NOR2BX1 U18679 ( .AN(n6944), .B(n7828), .Y(n6865) );
  XNOR2X1 U18680 ( .A(n6928), .B(n7800), .Y(n6748) );
  XNOR2X1 U18681 ( .A(n21054), .B(n25872), .Y(n6844) );
  OAI22X1 U18682 ( .A0(n6845), .A1(n6748), .B0(n6844), .B1(n6843), .Y(n6864)
         );
  XNOR2XL U18683 ( .A(n25869), .B(n25881), .Y(n6736) );
  XNOR2XL U18684 ( .A(n25869), .B(n7475), .Y(n6846) );
  OAI22XL U18685 ( .A0(n4592), .A1(n6736), .B0(n3046), .B1(n6846), .Y(n6863)
         );
  OAI22X1 U18686 ( .A0(n7093), .A1(n6734), .B0(n6780), .B1(n7094), .Y(n6743)
         );
  XNOR2X1 U18687 ( .A(n25867), .B(n25877), .Y(n6776) );
  OAI22X1 U18688 ( .A0(n6613), .A1(n6735), .B0(n7146), .B1(n6776), .Y(n6742)
         );
  OAI22XL U18689 ( .A0(n4592), .A1(n6737), .B0(n3046), .B1(n6736), .Y(n6741)
         );
  XOR2X1 U18690 ( .A(n6746), .B(M0_a_20_), .Y(n6745) );
  OAI22XL U18691 ( .A0(n4642), .A1(n7711), .B0(n7712), .B1(n6747), .Y(n6779)
         );
  OAI22XL U18692 ( .A0(n6845), .A1(n6749), .B0(n6748), .B1(n6843), .Y(n6790)
         );
  OAI22XL U18693 ( .A0(n6752), .A1(n7460), .B0(n7535), .B1(n6751), .Y(n6777)
         );
  OAI22X1 U18694 ( .A0(n7287), .A1(n6756), .B0(n6781), .B1(n7288), .Y(n6773)
         );
  XNOR2X1 U18695 ( .A(n23221), .B(n7164), .Y(n6774) );
  OAI22X1 U18696 ( .A0(n7633), .A1(n6757), .B0(n6774), .B1(n7634), .Y(n6772)
         );
  XNOR2X1 U18697 ( .A(n25868), .B(n25879), .Y(n6782) );
  OAI22XL U18698 ( .A0(n7511), .A1(n6758), .B0(n7512), .B1(n6782), .Y(n6771)
         );
  XNOR2X1 U18699 ( .A(n23221), .B(n25882), .Y(n6823) );
  OAI22XL U18700 ( .A0(n7633), .A1(n6774), .B0(n6823), .B1(n7634), .Y(n6868)
         );
  XNOR2X1 U18701 ( .A(n25867), .B(n25876), .Y(n6837) );
  OAI22XL U18702 ( .A0(n6613), .A1(n6776), .B0(n7146), .B1(n6837), .Y(n6866)
         );
  ADDFHX1 U18703 ( .A(n6779), .B(n4769), .CI(n6777), .CO(n6875), .S(n6762) );
  XNOR2XL U18704 ( .A(n7286), .B(n7621), .Y(n6822) );
  OAI22X1 U18705 ( .A0(n7287), .A1(n6781), .B0(n6822), .B1(n7288), .Y(n6817)
         );
  XNOR2X1 U18706 ( .A(n25868), .B(n7569), .Y(n6820) );
  OAI22XL U18707 ( .A0(n7511), .A1(n6782), .B0(n7512), .B1(n6820), .Y(n6816)
         );
  XNOR2XL U18708 ( .A(n23219), .B(n6944), .Y(n6783) );
  OAI22XL U18709 ( .A0(n6791), .A1(n7712), .B0(n4642), .B1(n6783), .Y(n6794)
         );
  XNOR2X1 U18710 ( .A(n25870), .B(n7165), .Y(n6824) );
  ADDHXL U18711 ( .A(n6789), .B(n6790), .CO(n6850), .S(n6778) );
  XNOR2XL U18712 ( .A(M0_b_2_), .B(n23219), .Y(n6848) );
  OAI22XL U18713 ( .A0(n6791), .A1(n4642), .B0(n6848), .B1(n7712), .Y(n6849)
         );
  ADDFHX1 U18714 ( .A(n6794), .B(n4756), .CI(n6792), .CO(n6882), .S(n6803) );
  XNOR2X1 U18715 ( .A(n23220), .B(n25879), .Y(n6862) );
  OAI22XL U18716 ( .A0(n7535), .A1(n6819), .B0(n6862), .B1(n7460), .Y(n6827)
         );
  XNOR2X1 U18717 ( .A(n25868), .B(n25878), .Y(n6832) );
  NAND2X4 U18718 ( .A(n7828), .B(n6821), .Y(n7829) );
  OAI22XL U18719 ( .A0(n7829), .A1(n6944), .B0(M0_b_1_), .B1(n7828), .Y(n6825)
         );
  XNOR2XL U18720 ( .A(n7286), .B(n25877), .Y(n6831) );
  OAI22XL U18721 ( .A0(n7287), .A1(n6822), .B0(n6831), .B1(n7288), .Y(n6840)
         );
  XNOR2X1 U18722 ( .A(n23221), .B(n25881), .Y(n6841) );
  XNOR2X1 U18723 ( .A(n25870), .B(n7164), .Y(n6842) );
  XNOR2XL U18724 ( .A(n25866), .B(n6828), .Y(n6921) );
  OAI22XL U18725 ( .A0(n6991), .A1(n6834), .B0(n6990), .B1(n6921), .Y(n6918)
         );
  XNOR2X1 U18726 ( .A(n3209), .B(n25874), .Y(n6833) );
  XNOR2XL U18727 ( .A(n3209), .B(M0_b_20_), .Y(n6919) );
  OAI22XL U18728 ( .A0(n6613), .A1(n6836), .B0(n7146), .B1(n6931), .Y(n6916)
         );
  XNOR2XL U18729 ( .A(n7286), .B(n6830), .Y(n6929) );
  XNOR2X1 U18730 ( .A(n25868), .B(n7621), .Y(n6920) );
  OAI22XL U18731 ( .A0(n7511), .A1(n6832), .B0(n7512), .B1(n6920), .Y(n6926)
         );
  XNOR2X1 U18732 ( .A(n23219), .B(n7165), .Y(n6930) );
  OAI22XL U18733 ( .A0(n6847), .A1(n4642), .B0(n6930), .B1(n7712), .Y(n6925)
         );
  OAI22XL U18734 ( .A0(n6991), .A1(n6835), .B0(n6990), .B1(n6834), .Y(n6870)
         );
  OAI22XL U18735 ( .A0(n6613), .A1(n6837), .B0(n7146), .B1(n6836), .Y(n6869)
         );
  XNOR2X1 U18736 ( .A(n23221), .B(n7475), .Y(n6941) );
  OAI22XL U18737 ( .A0(n7633), .A1(n6841), .B0(n6941), .B1(n6300), .Y(n6947)
         );
  XNOR2X1 U18738 ( .A(n25870), .B(n25882), .Y(n6923) );
  OAI22XL U18739 ( .A0(n7829), .A1(M0_b_1_), .B0(n7828), .B1(M0_b_2_), .Y(
        n6945) );
  OAI22XL U18740 ( .A0(n6845), .A1(n6844), .B0(n6843), .B1(n21054), .Y(n6859)
         );
  XNOR2XL U18741 ( .A(M0_b_9_), .B(n25869), .Y(n6858) );
  OAI22XL U18742 ( .A0(n6858), .A1(n3046), .B0(n4592), .B1(n6846), .Y(n6856)
         );
  OAI22XL U18743 ( .A0(n6848), .A1(n4642), .B0(n6847), .B1(n7712), .Y(n6855)
         );
  CMPR32X1 U18744 ( .A(n6851), .B(n6849), .C(n6850), .CO(n6885), .S(n6881) );
  CMPR32X1 U18745 ( .A(n6857), .B(n6856), .C(n6855), .CO(n6937), .S(n6886) );
  OAI22XL U18746 ( .A0(n6858), .A1(n4592), .B0(n3046), .B1(n6924), .Y(n6940)
         );
  OAI22XL U18747 ( .A0(n7535), .A1(n6862), .B0(n6922), .B1(n7460), .Y(n6942)
         );
  ADDFHX1 U18748 ( .A(n6868), .B(n6867), .CI(n6866), .CO(n6873), .S(n6876) );
  ADDFHX1 U18749 ( .A(n6870), .B(n6871), .CI(n6869), .CO(n6915), .S(n6872) );
  ADDFHX1 U18750 ( .A(n6874), .B(n6873), .CI(n6872), .CO(n6935), .S(n6892) );
  ADDFHX1 U18751 ( .A(n6883), .B(n6882), .CI(n6881), .CO(n6898), .S(n6894) );
  ADDFHX1 U18752 ( .A(n6889), .B(n6888), .CI(n6887), .CO(n6896), .S(n6904) );
  ADDFHX1 U18753 ( .A(n6892), .B(n6891), .CI(n6890), .CO(n6932), .S(n6901) );
  ADDFHX4 U18754 ( .A(n6898), .B(n6897), .CI(n6896), .CO(n6954), .S(n6899) );
  ADDFHX4 U18755 ( .A(n6904), .B(n6903), .CI(n6902), .CO(n6909), .S(n6908) );
  NAND2X2 U18756 ( .A(n6910), .B(n6909), .Y(n7021) );
  NAND2X2 U18757 ( .A(n6912), .B(n6911), .Y(n7014) );
  ADDFHX1 U18758 ( .A(n6915), .B(n6914), .CI(n6913), .CO(n6999), .S(n6951) );
  ADDFHX1 U18759 ( .A(n6918), .B(n6917), .CI(n6916), .CO(n6996), .S(n6949) );
  OAI22XL U18760 ( .A0(n7093), .A1(n6919), .B0(n6963), .B1(n7094), .Y(n6973)
         );
  XNOR2X1 U18761 ( .A(n25868), .B(n25877), .Y(n6964) );
  OAI22X1 U18762 ( .A0(n7511), .A1(n6920), .B0(n7512), .B1(n6964), .Y(n6972)
         );
  OAI22XL U18763 ( .A0(n6991), .A1(n6921), .B0(n6990), .B1(n25866), .Y(n6971)
         );
  XNOR2X1 U18764 ( .A(n23220), .B(n25878), .Y(n6967) );
  OAI22XL U18765 ( .A0(n7535), .A1(n6922), .B0(n6967), .B1(n7460), .Y(n6970)
         );
  XNOR2XL U18766 ( .A(n25869), .B(n25879), .Y(n6965) );
  OAI22XL U18767 ( .A0(n4592), .A1(n6924), .B0(n3046), .B1(n6965), .Y(n6968)
         );
  ADDFHX1 U18768 ( .A(n6926), .B(n6927), .CI(n6925), .CO(n6962), .S(n6948) );
  OAI22X1 U18769 ( .A0(n7829), .A1(M0_b_2_), .B0(n7828), .B1(n4806), .Y(n6993)
         );
  XNOR2X1 U18770 ( .A(n23219), .B(n7164), .Y(n6966) );
  OAI22XL U18771 ( .A0(n6613), .A1(n6931), .B0(n7146), .B1(n6978), .Y(n6974)
         );
  CMPR32X1 U18772 ( .A(n6944), .B(n6943), .C(n6942), .CO(n6986), .S(n6938) );
  ADDFHX1 U18773 ( .A(n6947), .B(n6946), .CI(n6945), .CO(n6985), .S(n6913) );
  ADDFHX4 U18774 ( .A(n6956), .B(n6954), .CI(n6955), .CO(n6957), .S(n6912) );
  NAND2X2 U18775 ( .A(n6958), .B(n6957), .Y(n7256) );
  NAND2XL U18776 ( .A(n5622), .B(n7256), .Y(n6959) );
  CMPR32X1 U18777 ( .A(n6962), .B(n6961), .C(n6960), .CO(n7132), .S(n6997) );
  XNOR2X1 U18778 ( .A(n25868), .B(n25876), .Y(n7051) );
  OAI22XL U18779 ( .A0(n4592), .A1(n6965), .B0(n3046), .B1(n7028), .Y(n7032)
         );
  XNOR2X1 U18780 ( .A(n23219), .B(n25882), .Y(n7025) );
  OAI22X2 U18781 ( .A0(n4642), .A1(n6966), .B0(n7025), .B1(n7712), .Y(n7036)
         );
  XNOR2X1 U18782 ( .A(n23220), .B(n7621), .Y(n7038) );
  OAI22XL U18783 ( .A0(n7535), .A1(n6967), .B0(n7038), .B1(n7460), .Y(n7035)
         );
  ADDFHX1 U18784 ( .A(n6970), .B(n6969), .CI(n6968), .CO(n7075), .S(n6994) );
  XNOR2XL U18785 ( .A(n7286), .B(M0_b_18_), .Y(n7024) );
  OAI22XL U18786 ( .A0(n7287), .A1(n6976), .B0(n7024), .B1(n7288), .Y(n7031)
         );
  OAI22XL U18787 ( .A0(n6613), .A1(n6978), .B0(n7146), .B1(n7039), .Y(n7029)
         );
  INVXL U18788 ( .A(n7257), .Y(n7005) );
  NOR2XL U18789 ( .A(n7009), .B(n7020), .Y(n7012) );
  OAI21XL U18790 ( .A0(n7010), .A1(n7020), .B0(n7021), .Y(n7011) );
  OAI22XL U18791 ( .A0(n7287), .A1(n7024), .B0(n7065), .B1(n7288), .Y(n7064)
         );
  XNOR2X1 U18792 ( .A(n23219), .B(n25881), .Y(n7047) );
  XNOR2X1 U18793 ( .A(n23221), .B(n25879), .Y(n7061) );
  OAI22XL U18794 ( .A0(n7633), .A1(n7026), .B0(n7061), .B1(n7634), .Y(n7062)
         );
  OAI22X1 U18795 ( .A0(n7829), .A1(n7165), .B0(n7828), .B1(n7164), .Y(n7045)
         );
  OAI22XL U18796 ( .A0(n4592), .A1(n7028), .B0(n3046), .B1(n7066), .Y(n7044)
         );
  ADDFHX1 U18797 ( .A(n7034), .B(n7033), .CI(n7032), .CO(n7086), .S(n7073) );
  XNOR2X1 U18798 ( .A(n25867), .B(n7800), .Y(n7048) );
  OAI22X1 U18799 ( .A0(n6613), .A1(n7039), .B0(n7146), .B1(n7048), .Y(n7042)
         );
  OAI2BB1XL U18800 ( .A0N(n7040), .A1N(n6991), .B0(n25866), .Y(n7041) );
  ADDFHX1 U18801 ( .A(n7043), .B(n7042), .CI(n7041), .CO(n7110), .S(n7084) );
  XNOR2X1 U18802 ( .A(n23219), .B(n7475), .Y(n7114) );
  OAI22XL U18803 ( .A0(n4642), .A1(n7047), .B0(n7114), .B1(n7712), .Y(n7113)
         );
  XNOR2X1 U18804 ( .A(n25868), .B(n7646), .Y(n7050) );
  XNOR2X1 U18805 ( .A(n25868), .B(n25875), .Y(n7091) );
  OAI22XL U18806 ( .A0(n6613), .A1(n7048), .B0(n7146), .B1(n7088), .Y(n7111)
         );
  XNOR2X1 U18807 ( .A(n23220), .B(n25876), .Y(n7095) );
  OAI22XL U18808 ( .A0(n7535), .A1(n7049), .B0(n7095), .B1(n7460), .Y(n7117)
         );
  XNOR2XL U18809 ( .A(M0_b_9_), .B(n25870), .Y(n7053) );
  XNOR2X1 U18810 ( .A(n25870), .B(n25880), .Y(n7089) );
  CMPR32X1 U18811 ( .A(n4806), .B(M0_b_2_), .C(n7054), .CO(n7115), .S(n7068)
         );
  NAND2BXL U18812 ( .AN(n7057), .B(n7056), .Y(n7060) );
  XNOR2X1 U18813 ( .A(n23221), .B(n7569), .Y(n7090) );
  XNOR2XL U18814 ( .A(n7286), .B(n25873), .Y(n7087) );
  OAI22XL U18815 ( .A0(n7287), .A1(n7065), .B0(n7087), .B1(n7288), .Y(n7101)
         );
  ADDFHX1 U18816 ( .A(n7069), .B(n7068), .CI(n7067), .CO(n7103), .S(n7129) );
  CMPR32X1 U18817 ( .A(n7086), .B(n7085), .C(n7084), .CO(n7119), .S(n7240) );
  XNOR2X1 U18818 ( .A(n7286), .B(n7800), .Y(n7166) );
  OAI22XL U18819 ( .A0(n7287), .A1(n7087), .B0(n7166), .B1(n7288), .Y(n7158)
         );
  XNOR2X1 U18820 ( .A(n23221), .B(n25878), .Y(n7167) );
  OAI22XL U18821 ( .A0(n7633), .A1(n7090), .B0(n7167), .B1(n7634), .Y(n7144)
         );
  XNOR2X1 U18822 ( .A(n25868), .B(n25874), .Y(n7147) );
  OAI22XL U18823 ( .A0(n7511), .A1(n7091), .B0(n7512), .B1(n7147), .Y(n7143)
         );
  OAI2BB1XL U18824 ( .A0N(n7094), .A1N(n7093), .B0(n7092), .Y(n7142) );
  XNOR2X1 U18825 ( .A(n23220), .B(n7646), .Y(n7145) );
  OAI22XL U18826 ( .A0(n7535), .A1(n7095), .B0(n7145), .B1(n7460), .Y(n7163)
         );
  ADDFHX1 U18827 ( .A(n7107), .B(n7106), .CI(n7105), .CO(n7170), .S(n7102) );
  CMPR32X1 U18828 ( .A(n7110), .B(n7109), .C(n7108), .CO(n7169), .S(n7118) );
  OAI22XL U18829 ( .A0(n7829), .A1(n25882), .B0(n7828), .B1(n25881), .Y(n7161)
         );
  XNOR2XL U18830 ( .A(M0_b_9_), .B(n23219), .Y(n7162) );
  OAI22XL U18831 ( .A0(n7162), .A1(n7712), .B0(n4642), .B1(n7114), .Y(n7159)
         );
  ADDFHX1 U18832 ( .A(n7117), .B(n7116), .CI(n7115), .CO(n7139), .S(n7104) );
  CMPR32X1 U18833 ( .A(n7129), .B(n7128), .C(n7127), .CO(n7122), .S(n7247) );
  CMPR32X1 U18834 ( .A(n7132), .B(n7131), .C(n7130), .CO(n7246), .S(n7254) );
  NOR2X2 U18835 ( .A(n7263), .B(n7262), .Y(n7317) );
  CMPR32X1 U18836 ( .A(n7138), .B(n7137), .C(n7136), .CO(n7173), .S(n7153) );
  OAI22X2 U18837 ( .A0(n6613), .A1(n25867), .B0(n7146), .B1(n6829), .Y(n7195)
         );
  XNOR2X1 U18838 ( .A(n25868), .B(n25873), .Y(n7189) );
  OAI22XL U18839 ( .A0(n7511), .A1(n7147), .B0(n7512), .B1(n7189), .Y(n7194)
         );
  OAI22XL U18840 ( .A0(n7829), .A1(n25881), .B0(n7828), .B1(n7475), .Y(n7182)
         );
  OAI22XL U18841 ( .A0(n4592), .A1(n7149), .B0(n3046), .B1(n7185), .Y(n7180)
         );
  CMPR32X1 U18842 ( .A(n7155), .B(n7154), .C(n7153), .CO(n7176), .S(n7152) );
  XNOR2X1 U18843 ( .A(n23219), .B(n25880), .Y(n7183) );
  OAI22XL U18844 ( .A0(n7162), .A1(n4642), .B0(n7183), .B1(n7712), .Y(n7188)
         );
  CMPR32X1 U18845 ( .A(n7165), .B(n7164), .C(n7163), .CO(n7187), .S(n7138) );
  INVXL U18846 ( .A(n25882), .Y(n7193) );
  XNOR2X1 U18847 ( .A(n7286), .B(n25872), .Y(n7190) );
  OAI22XL U18848 ( .A0(n7633), .A1(n7167), .B0(n7197), .B1(n6300), .Y(n7191)
         );
  ADDFHX1 U18849 ( .A(n7182), .B(n7181), .CI(n7180), .CO(n7215), .S(n7198) );
  XNOR2X1 U18850 ( .A(n23219), .B(n25879), .Y(n7226) );
  OAI22XL U18851 ( .A0(n4642), .A1(n7183), .B0(n7226), .B1(n7712), .Y(n7218)
         );
  OAI22XL U18852 ( .A0(n4592), .A1(n7185), .B0(n3046), .B1(n7222), .Y(n7216)
         );
  XNOR2X1 U18853 ( .A(n25868), .B(n7800), .Y(n7221) );
  OAI22XL U18854 ( .A0(n7511), .A1(n7189), .B0(n7512), .B1(n7221), .Y(n7224)
         );
  OAI22XL U18855 ( .A0(n7287), .A1(n7190), .B0(n7288), .B1(n4789), .Y(n7231)
         );
  ADDFHX1 U18856 ( .A(n7193), .B(n7192), .CI(n7191), .CO(n7230), .S(n7186) );
  ADDFHX4 U18857 ( .A(n7196), .B(n7195), .CI(n7194), .CO(n7229), .S(n7199) );
  OAI22X1 U18858 ( .A0(n7829), .A1(n7475), .B0(M0_b_9_), .B1(n7828), .Y(n7234)
         );
  NOR2X2 U18859 ( .A(n7267), .B(n7266), .Y(n7447) );
  ADDFHX1 U18860 ( .A(n7206), .B(n7205), .CI(n7204), .CO(n7269), .S(n7267) );
  CMPR32X1 U18861 ( .A(n7215), .B(n7214), .C(n7213), .CO(n7279), .S(n7211) );
  ADDFHX1 U18862 ( .A(n7218), .B(n7217), .CI(n7216), .CO(n7282), .S(n7214) );
  XNOR2X1 U18863 ( .A(n23220), .B(n25873), .Y(n7291) );
  OAI22XL U18864 ( .A0(n7535), .A1(n7219), .B0(n7291), .B1(n7460), .Y(n7285)
         );
  XNOR2X1 U18865 ( .A(n25868), .B(n25872), .Y(n7289) );
  XNOR2XL U18866 ( .A(n25869), .B(n25875), .Y(n7293) );
  OAI22XL U18867 ( .A0(n4592), .A1(n7222), .B0(n3046), .B1(n7293), .Y(n7283)
         );
  CMPR32X1 U18868 ( .A(n7225), .B(n7224), .C(n7223), .CO(n7280), .S(n7209) );
  XNOR2X1 U18869 ( .A(n23219), .B(n7569), .Y(n7297) );
  OAI22XL U18870 ( .A0(n4642), .A1(n7226), .B0(n7297), .B1(n7712), .Y(n7296)
         );
  OAI22XL U18871 ( .A0(n7829), .A1(M0_b_9_), .B0(n7828), .B1(n25880), .Y(n7295) );
  INVXL U18872 ( .A(n7475), .Y(n7300) );
  OAI22XL U18873 ( .A0(n7287), .A1(n4789), .B0(n7288), .B1(n3213), .Y(n7299)
         );
  OAI22XL U18874 ( .A0(n7633), .A1(n7232), .B0(n7290), .B1(n6300), .Y(n7298)
         );
  ADDFHX2 U18875 ( .A(n7245), .B(n7244), .CI(n7243), .CO(n7250), .S(n7252) );
  CMPR32X1 U18876 ( .A(n7248), .B(n7247), .C(n7246), .CO(n7237), .S(n7249) );
  ADDFHX1 U18877 ( .A(n7273), .B(n7272), .CI(n7271), .CO(n7305), .S(n7268) );
  CMPR32X1 U18878 ( .A(n7276), .B(n7275), .C(n7274), .CO(n7455), .S(n7277) );
  CMPR32X1 U18879 ( .A(n7282), .B(n7281), .C(n7280), .CO(n7481), .S(n7278) );
  OAI2BB1XL U18880 ( .A0N(n7288), .A1N(n7287), .B0(n7286), .Y(n7473) );
  OAI22XL U18881 ( .A0(n7511), .A1(n7289), .B0(n7512), .B1(n25868), .Y(n7472)
         );
  OAI22XL U18882 ( .A0(n7633), .A1(n7290), .B0(n7459), .B1(n6300), .Y(n7471)
         );
  XNOR2X1 U18883 ( .A(n23220), .B(n7800), .Y(n7461) );
  XNOR2X1 U18884 ( .A(n25870), .B(n25877), .Y(n7467) );
  OAI22XL U18885 ( .A0(n4592), .A1(n7293), .B0(n3046), .B1(n7466), .Y(n7462)
         );
  OAI22XL U18886 ( .A0(n7829), .A1(n25880), .B0(n7828), .B1(n25879), .Y(n7478)
         );
  XNOR2X1 U18887 ( .A(n23219), .B(n25878), .Y(n7465) );
  INVXL U18888 ( .A(n7487), .Y(n7306) );
  INVXL U18889 ( .A(n7324), .Y(n7309) );
  INVXL U18890 ( .A(n7312), .Y(n7314) );
  NAND2XL U18891 ( .A(n7314), .B(n7313), .Y(n7315) );
  XNOR2X1 U18892 ( .A(n7316), .B(n7315), .Y(n10737) );
  INVXL U18893 ( .A(n7320), .Y(n7323) );
  NAND2XL U18894 ( .A(n7325), .B(n7324), .Y(n7326) );
  OAI21XL U18895 ( .A0(n7352), .A1(n7353), .B0(n7355), .Y(n7328) );
  OAI21XL U18896 ( .A0(M0_U4_U1_enc_tree_2__4__16_), .A1(
        M0_U3_U1_enc_tree_2__4__16_), .B0(n7328), .Y(n7337) );
  INVXL U18897 ( .A(n7360), .Y(n7363) );
  INVXL U18898 ( .A(n7361), .Y(n7362) );
  INVXL U18899 ( .A(n7365), .Y(n7367) );
  NAND2XL U18900 ( .A(n7367), .B(n7366), .Y(n7368) );
  OAI21XL U18901 ( .A0(n6266), .A1(n26290), .B0(n24022), .Y(n7371) );
  NOR2X1 U18902 ( .A(n7371), .B(n7370), .Y(n7843) );
  OAI21XL U18903 ( .A0(n6266), .A1(n26291), .B0(n14407), .Y(n7373) );
  OR2X2 U18904 ( .A(n7843), .B(n7842), .Y(n7399) );
  OAI21XL U18905 ( .A0(n6266), .A1(n26289), .B0(n25216), .Y(n7375) );
  OAI21XL U18906 ( .A0(n6266), .A1(n26299), .B0(n25213), .Y(n7379) );
  OAI21XL U18907 ( .A0(n6266), .A1(n26305), .B0(n25210), .Y(n7384) );
  NOR2X1 U18908 ( .A(n7384), .B(n7383), .Y(n7849) );
  AOI2BB2X1 U18909 ( .B0(n7868), .B1(n7869), .A0N(n7869), .A1N(n7868), .Y(
        n10721) );
  CMPR32X1 U18910 ( .A(n7853), .B(n7403), .C(n7402), .CO(n7868), .S(n23685) );
  CMPR32X1 U18911 ( .A(n7857), .B(n7407), .C(n7406), .CO(n7414), .S(n23822) );
  CMPR32X1 U18912 ( .A(n7859), .B(n7409), .C(n7408), .CO(n7410), .S(n23865) );
  CMPR32X1 U18913 ( .A(n7856), .B(n7411), .C(n7410), .CO(n7406), .S(n23782) );
  CMPR22X1 U18914 ( .A(n7843), .B(n7858), .CO(n7408), .S(n23862) );
  CMPR32X1 U18915 ( .A(n7855), .B(n7413), .C(n7412), .CO(n7404), .S(n23683) );
  CMPR32X1 U18916 ( .A(n7854), .B(n7415), .C(n7414), .CO(n7412), .S(n23854) );
  NAND4BXL U18917 ( .AN(n23850), .B(n7418), .C(n7417), .D(n7416), .Y(n7419) );
  INVXL U18918 ( .A(n7872), .Y(n7421) );
  NAND2XL U18919 ( .A(n7426), .B(n7442), .Y(n7428) );
  INVXL U18920 ( .A(n7424), .Y(n7425) );
  INVXL U18921 ( .A(n7429), .Y(n7431) );
  NOR2XL U18922 ( .A(n3168), .B(n7447), .Y(n7435) );
  INVXL U18923 ( .A(n7444), .Y(n7433) );
  OAI21XL U18924 ( .A0(n7433), .A1(n7447), .B0(n7448), .Y(n7434) );
  INVXL U18925 ( .A(n7438), .Y(n7440) );
  INVXL U18926 ( .A(n7447), .Y(n7449) );
  ADDFHX1 U18927 ( .A(n7455), .B(n7454), .CI(n7453), .CO(n7483), .S(n7304) );
  ADDFHX1 U18928 ( .A(n7458), .B(n7457), .CI(n7456), .CO(n7493), .S(n7479) );
  INVXL U18929 ( .A(n25880), .Y(n7500) );
  XNOR2X1 U18930 ( .A(n23220), .B(n25872), .Y(n7509) );
  OAI22XL U18931 ( .A0(n7535), .A1(n7461), .B0(n7509), .B1(n7460), .Y(n7498)
         );
  XNOR2X1 U18932 ( .A(n23219), .B(n7621), .Y(n7507) );
  OAI22XL U18933 ( .A0(n4642), .A1(n7465), .B0(n7507), .B1(n7712), .Y(n7503)
         );
  XNOR2XL U18934 ( .A(n25869), .B(n25873), .Y(n7510) );
  ADDFHX1 U18935 ( .A(n7470), .B(n7469), .CI(n7468), .CO(n7517), .S(n7480) );
  OAI22XL U18936 ( .A0(n7829), .A1(n25879), .B0(n7828), .B1(n7569), .Y(n7515)
         );
  OAI22XL U18937 ( .A0(n7511), .A1(n25868), .B0(n7512), .B1(n6476), .Y(n7514)
         );
  CMPR32X1 U18938 ( .A(n7475), .B(M0_b_9_), .C(n7474), .CO(n7513), .S(n7477)
         );
  CMPR32X1 U18939 ( .A(n7481), .B(n7480), .C(n7479), .CO(n7491), .S(n7453) );
  NOR2X1 U18940 ( .A(n7483), .B(n7482), .Y(n7490) );
  INVXL U18941 ( .A(n7490), .Y(n7484) );
  INVXL U18942 ( .A(n7779), .Y(n7753) );
  ADDFHX2 U18943 ( .A(n7496), .B(n7495), .CI(n7494), .CO(n7610), .S(n7516) );
  OAI22XL U18944 ( .A0(n7633), .A1(n7497), .B0(n7536), .B1(n6300), .Y(n7533)
         );
  ADDFHX1 U18945 ( .A(n7500), .B(n7499), .CI(n7498), .CO(n7538), .S(n7506) );
  ADDFHX1 U18946 ( .A(n7503), .B(n7502), .CI(n7501), .CO(n7537), .S(n7504) );
  ADDFHX4 U18947 ( .A(n7506), .B(n7505), .CI(n7504), .CO(n7597), .S(n7518) );
  OAI22XL U18948 ( .A0(n4642), .A1(n7507), .B0(n7530), .B1(n7712), .Y(n7529)
         );
  OAI22XL U18949 ( .A0(n7535), .A1(n7509), .B0(n7556), .B1(n23220), .Y(n7526)
         );
  OAI2BB1XL U18950 ( .A0N(n7512), .A1N(n7511), .B0(n25868), .Y(n7524) );
  CMPR32X1 U18951 ( .A(n7515), .B(n7514), .C(n7513), .CO(n7540), .S(n7495) );
  NOR2XL U18952 ( .A(n7520), .B(n7521), .Y(n7519) );
  NAND2X1 U18953 ( .A(n7521), .B(n7520), .Y(n7657) );
  XNOR2X2 U18954 ( .A(n7523), .B(n7522), .Y(n20830) );
  ADDFHX1 U18955 ( .A(n7526), .B(n7525), .CI(n7524), .CO(n7595), .S(n7541) );
  ADDFHX1 U18956 ( .A(n7529), .B(n7528), .CI(n7527), .CO(n7594), .S(n7542) );
  XNOR2X1 U18957 ( .A(n23219), .B(n25876), .Y(n7554) );
  OAI22XL U18958 ( .A0(n4642), .A1(n7530), .B0(n7554), .B1(n7712), .Y(n7553)
         );
  OAI22XL U18959 ( .A0(n7829), .A1(n25878), .B0(n7828), .B1(n7621), .Y(n7545)
         );
  CMPR32X1 U18960 ( .A(n25879), .B(n25880), .C(n7533), .CO(n7544), .S(n7539)
         );
  OAI22XL U18961 ( .A0(n7535), .A1(n23220), .B0(n7460), .B1(n7534), .Y(n7549)
         );
  OAI22XL U18962 ( .A0(n7633), .A1(n7536), .B0(n7547), .B1(n6300), .Y(n7548)
         );
  ADDFHX1 U18963 ( .A(n7539), .B(n7538), .CI(n7537), .CO(n7600), .S(n7598) );
  ADDFHX1 U18964 ( .A(n7542), .B(n7541), .CI(n7540), .CO(n7599), .S(n7596) );
  ADDFHX1 U18965 ( .A(n7545), .B(n7544), .CI(n7543), .CO(n7562), .S(n7601) );
  OAI22XL U18966 ( .A0(n7829), .A1(n7621), .B0(n7828), .B1(n25877), .Y(n7567)
         );
  OAI22XL U18967 ( .A0(n7633), .A1(n7547), .B0(n7570), .B1(n6300), .Y(n7568)
         );
  CMPR32X1 U18968 ( .A(n7553), .B(n7552), .C(n7551), .CO(n7558), .S(n7593) );
  XNOR2X1 U18969 ( .A(n23219), .B(n7646), .Y(n7571) );
  OAI22XL U18970 ( .A0(n4642), .A1(n7554), .B0(n7571), .B1(n7712), .Y(n7574)
         );
  OAI2BB1XL U18971 ( .A0N(n7556), .A1N(n7535), .B0(n23220), .Y(n7572) );
  CMPR32X1 U18972 ( .A(n7562), .B(n7561), .C(n7560), .CO(n7576), .S(n7602) );
  OAI22XL U18973 ( .A0(n7829), .A1(n25877), .B0(n7828), .B1(n25876), .Y(n7586)
         );
  OAI22XL U18974 ( .A0(n4592), .A1(n25869), .B0(n3046), .B1(n7564), .Y(n7584)
         );
  CMPR32X1 U18975 ( .A(n7567), .B(n7566), .C(n7565), .CO(n7582), .S(n7561) );
  CMPR32X1 U18976 ( .A(n7569), .B(n25878), .C(n7568), .CO(n7580), .S(n7565) );
  OAI22XL U18977 ( .A0(n4642), .A1(n7571), .B0(n7587), .B1(n7712), .Y(n7590)
         );
  ADDFHX1 U18978 ( .A(n7580), .B(n7579), .CI(n7578), .CO(n7653), .S(n7581) );
  XNOR2X1 U18979 ( .A(n23219), .B(n25874), .Y(n7616) );
  OAI22XL U18980 ( .A0(n4642), .A1(n7587), .B0(n7616), .B1(n7712), .Y(n7619)
         );
  OAI2BB1XL U18981 ( .A0N(n3046), .A1N(n4592), .B0(M0_a_15_), .Y(n7617) );
  OAI22XL U18982 ( .A0(n7633), .A1(n7589), .B0(n7634), .B1(n23221), .Y(n7620)
         );
  NOR2X2 U18983 ( .A(n7666), .B(n7665), .Y(n7768) );
  CMPR32X1 U18984 ( .A(n7604), .B(n7603), .C(n7602), .CO(n7664), .S(n7661) );
  OR2X2 U18985 ( .A(n7662), .B(n7661), .Y(n7786) );
  CMPR32X1 U18986 ( .A(n7607), .B(n7606), .C(n7605), .CO(n7662), .S(n7659) );
  CMPR32X1 U18987 ( .A(n7610), .B(n7609), .C(n7608), .CO(n7658), .S(n7521) );
  NAND2X1 U18988 ( .A(n7776), .B(n7772), .Y(n7752) );
  XNOR2X1 U18989 ( .A(n23219), .B(n25873), .Y(n7628) );
  OAI22XL U18990 ( .A0(n4642), .A1(n7616), .B0(n7628), .B1(n7712), .Y(n7629)
         );
  CMPR32X1 U18991 ( .A(n7619), .B(n7618), .C(n7617), .CO(n7636), .S(n7623) );
  OAI22XL U18992 ( .A0(n7829), .A1(n7646), .B0(n7828), .B1(n25875), .Y(n7627)
         );
  CMPR32X1 U18993 ( .A(n25877), .B(n7621), .C(n7620), .CO(n7625), .S(n7613) );
  CMPR32X1 U18994 ( .A(n7627), .B(n7626), .C(n7625), .CO(n7640), .S(n7635) );
  XNOR2X1 U18995 ( .A(n23219), .B(n7800), .Y(n7647) );
  OAI22XL U18996 ( .A0(n4642), .A1(n7628), .B0(n7647), .B1(n7712), .Y(n7645)
         );
  OR2X2 U18997 ( .A(n7676), .B(n7675), .Y(n7807) );
  CMPR32X1 U18998 ( .A(n25876), .B(n7646), .C(n7645), .CO(n7693), .S(n7650) );
  XNOR2X1 U18999 ( .A(n23219), .B(n25872), .Y(n7696) );
  OAI22XL U19000 ( .A0(n7829), .A1(n25874), .B0(n7828), .B1(n25873), .Y(n7689)
         );
  CMPR32X1 U19001 ( .A(n7650), .B(n7649), .C(n7648), .CO(n7686), .S(n7639) );
  CMPR32X1 U19002 ( .A(n7653), .B(n7652), .C(n7651), .CO(n7674), .S(n7665) );
  CMPR32X1 U19003 ( .A(n7656), .B(n7655), .C(n7654), .CO(n7676), .S(n7673) );
  INVXL U19004 ( .A(n7722), .Y(n7683) );
  NOR2XL U19005 ( .A(n7815), .B(n7683), .Y(n7701) );
  INVXL U19006 ( .A(n7701), .Y(n7685) );
  NAND2XL U19007 ( .A(n7659), .B(n7658), .Y(n7775) );
  INVXL U19008 ( .A(n7775), .Y(n7660) );
  AOI21X1 U19009 ( .A0(n7776), .A1(n7771), .B0(n7660), .Y(n7754) );
  NAND2XL U19010 ( .A(n7662), .B(n7661), .Y(n7785) );
  INVXL U19011 ( .A(n7785), .Y(n7755) );
  NAND2XL U19012 ( .A(n7666), .B(n7665), .Y(n7769) );
  OAI21XL U19013 ( .A0(n7768), .A1(n7762), .B0(n7769), .Y(n7667) );
  NAND2XL U19014 ( .A(n7678), .B(n7677), .Y(n7811) );
  INVXL U19015 ( .A(n7811), .Y(n7679) );
  INVXL U19016 ( .A(n7728), .Y(n7682) );
  INVXL U19017 ( .A(n7704), .Y(n7684) );
  CMPR32X1 U19018 ( .A(n7688), .B(n7687), .C(n7686), .CO(n7698), .S(n7677) );
  CMPR32X1 U19019 ( .A(n7694), .B(n7693), .C(n7692), .CO(n7708), .S(n7687) );
  NAND2XL U19020 ( .A(n7701), .B(n7703), .Y(n7706) );
  CMPR32X1 U19021 ( .A(n7709), .B(n7708), .C(n7707), .CO(n7717), .S(n7697) );
  CMPR32X1 U19022 ( .A(n25874), .B(n25875), .C(n7710), .CO(n7735), .S(n7713)
         );
  CMPR32X1 U19023 ( .A(n7715), .B(n7714), .C(n7713), .CO(n7733), .S(n7707) );
  INVXL U19024 ( .A(n7815), .Y(n7789) );
  INVXL U19025 ( .A(n7788), .Y(n7730) );
  NAND2XL U19026 ( .A(n7789), .B(n7730), .Y(n7732) );
  OAI21XL U19027 ( .A0(n7725), .A1(n7724), .B0(n7723), .Y(n7726) );
  INVXL U19028 ( .A(n7792), .Y(n7729) );
  AOI21X1 U19029 ( .A0(n7793), .A1(n7730), .B0(n7729), .Y(n7731) );
  OAI21X1 U19030 ( .A0(n3494), .A1(n7732), .B0(n7731), .Y(n7743) );
  CMPR32X1 U19031 ( .A(n7735), .B(n7734), .C(n7733), .CO(n7740), .S(n7716) );
  OAI2BB1X1 U19032 ( .A0N(n7712), .A1N(n4642), .B0(n23219), .Y(n7798) );
  CMPR32X1 U19033 ( .A(n7738), .B(n7737), .C(n7736), .CO(n7796), .S(n7734) );
  XNOR2X2 U19034 ( .A(n7743), .B(n7742), .Y(n20372) );
  INVXL U19035 ( .A(n7805), .Y(n7748) );
  OAI21X1 U19036 ( .A0(n7822), .A1(n7746), .B0(n7745), .Y(n7808) );
  INVXL U19037 ( .A(n7808), .Y(n7747) );
  INVXL U19038 ( .A(n7752), .Y(n7781) );
  NAND2XL U19039 ( .A(n7781), .B(n7786), .Y(n7758) );
  NOR2XL U19040 ( .A(n7753), .B(n7758), .Y(n7761) );
  INVXL U19041 ( .A(n7761), .Y(n7760) );
  INVXL U19042 ( .A(n7754), .Y(n7780) );
  AOI21XL U19043 ( .A0(n7780), .A1(n7786), .B0(n7755), .Y(n7756) );
  OAI21XL U19044 ( .A0(n7758), .A1(n7757), .B0(n7756), .Y(n7765) );
  INVXL U19045 ( .A(n7765), .Y(n7759) );
  NAND2XL U19046 ( .A(n7761), .B(n7764), .Y(n7767) );
  INVXL U19047 ( .A(n7762), .Y(n7763) );
  AOI21XL U19048 ( .A0(n7765), .A1(n7764), .B0(n7763), .Y(n7766) );
  NAND2XL U19049 ( .A(n7779), .B(n7772), .Y(n7774) );
  AOI21XL U19050 ( .A0(n7782), .A1(n7772), .B0(n7771), .Y(n7773) );
  XNOR2X2 U19051 ( .A(n7778), .B(n7777), .Y(n20832) );
  NAND2XL U19052 ( .A(n7779), .B(n7781), .Y(n7784) );
  AOI21XL U19053 ( .A0(n7782), .A1(n7781), .B0(n7780), .Y(n7783) );
  OAI21X1 U19054 ( .A0(n3605), .A1(n7784), .B0(n7783), .Y(n7787) );
  NAND2XL U19055 ( .A(n7789), .B(n7814), .Y(n7795) );
  AOI21XL U19056 ( .A0(n7793), .A1(n7814), .B0(n7819), .Y(n7794) );
  CMPR32X1 U19057 ( .A(n7798), .B(n7797), .C(n7796), .CO(n7802), .S(n7739) );
  CMPR32X1 U19058 ( .A(n25873), .B(n7800), .C(n7799), .CO(n7825), .S(n7797) );
  OR2X2 U19059 ( .A(n7802), .B(n7801), .Y(n7818) );
  CMPR32X1 U19060 ( .A(n7827), .B(n7826), .C(n7825), .CO(n7832), .S(n7801) );
  INVXL U19061 ( .A(n10721), .Y(n7867) );
  NAND3XL U19062 ( .A(n7844), .B(n7843), .C(n7842), .Y(n7866) );
  OAI21XL U19063 ( .A0(n7866), .A1(n7865), .B0(n7864), .Y(n23198) );
  AOI21XL U19064 ( .A0(n23683), .A1(n23864), .B0(n23863), .Y(n7879) );
  NOR2XL U19065 ( .A(n25886), .B(cs[1]), .Y(n23072) );
  NOR2X4 U19066 ( .A(n25887), .B(cs[0]), .Y(n7885) );
  INVX8 U19067 ( .A(n21111), .Y(n19161) );
  AOI22XL U19068 ( .A0(y10[30]), .A1(n19235), .B0(n19161), .B1(temp1[30]), .Y(
        n7883) );
  INVXL U19069 ( .A(n8192), .Y(n7890) );
  NAND2X2 U19070 ( .A(n7885), .B(n25886), .Y(n24632) );
  NAND2X1 U19071 ( .A(n7890), .B(n8148), .Y(n23690) );
  NAND2XL U19072 ( .A(n6217), .B(y10[3]), .Y(n7894) );
  NAND2XL U19073 ( .A(n19216), .B(w1[35]), .Y(n7892) );
  NAND2XL U19074 ( .A(n3120), .B(y20[3]), .Y(n7891) );
  AOI22XL U19075 ( .A0(n19346), .A1(y10[3]), .B0(n3062), .B1(temp1[3]), .Y(
        n7895) );
  OAI21XL U19076 ( .A0(n3063), .A1(n26590), .B0(n7895), .Y(n8424) );
  NOR2XL U19077 ( .A(n8459), .B(n8424), .Y(n7917) );
  NAND2XL U19078 ( .A(n6217), .B(y10[2]), .Y(n7899) );
  NAND2XL U19079 ( .A(n19216), .B(w1[34]), .Y(n7897) );
  NAND2XL U19080 ( .A(n3120), .B(y20[2]), .Y(n7896) );
  AOI22XL U19081 ( .A0(n19346), .A1(y10[2]), .B0(n3062), .B1(temp1[2]), .Y(
        n7900) );
  OAI21XL U19082 ( .A0(n3063), .A1(n26591), .B0(n7900), .Y(n8422) );
  NOR2XL U19083 ( .A(n8443), .B(n8422), .Y(n7901) );
  NOR2XL U19084 ( .A(n7917), .B(n7901), .Y(n7920) );
  NAND2XL U19085 ( .A(n19216), .B(w1[33]), .Y(n7903) );
  NAND2XL U19086 ( .A(n3120), .B(y20[1]), .Y(n7902) );
  AOI22XL U19087 ( .A0(n19349), .A1(y10[1]), .B0(n3026), .B1(temp1[1]), .Y(
        n7906) );
  OAI21XL U19088 ( .A0(n3063), .A1(n26592), .B0(n7906), .Y(n8479) );
  NOR2XL U19089 ( .A(n8509), .B(n8479), .Y(n7914) );
  NAND2XL U19090 ( .A(n6217), .B(y10[0]), .Y(n7910) );
  NAND2XL U19091 ( .A(n3027), .B(w2[0]), .Y(n7909) );
  NAND2XL U19092 ( .A(n19216), .B(w1[32]), .Y(n7908) );
  NAND2XL U19093 ( .A(n3120), .B(y20[0]), .Y(n7907) );
  AOI22XL U19094 ( .A0(n19346), .A1(y10[0]), .B0(n19216), .B1(temp1[0]), .Y(
        n7911) );
  OAI21XL U19095 ( .A0(n3063), .A1(n26593), .B0(n7911), .Y(n8477) );
  NAND2XL U19096 ( .A(n8496), .B(n8477), .Y(n7913) );
  NAND2XL U19097 ( .A(n8509), .B(n8479), .Y(n7912) );
  OAI21XL U19098 ( .A0(n7914), .A1(n7913), .B0(n7912), .Y(n7919) );
  NAND2XL U19099 ( .A(n8443), .B(n8422), .Y(n7916) );
  NAND2XL U19100 ( .A(n8459), .B(n8424), .Y(n7915) );
  OAI21XL U19101 ( .A0(n7917), .A1(n7916), .B0(n7915), .Y(n7918) );
  NAND2XL U19102 ( .A(n6217), .B(y10[4]), .Y(n7924) );
  NAND2XL U19103 ( .A(n3062), .B(w1[36]), .Y(n7922) );
  NAND2XL U19104 ( .A(n3120), .B(y20[4]), .Y(n7921) );
  AOI22XL U19105 ( .A0(n19346), .A1(y10[4]), .B0(n3026), .B1(temp1[4]), .Y(
        n7925) );
  OAI21XL U19106 ( .A0(n19237), .A1(n26589), .B0(n7925), .Y(n8427) );
  NOR2XL U19107 ( .A(n8474), .B(n8427), .Y(n7931) );
  NAND2XL U19108 ( .A(n6217), .B(y10[5]), .Y(n7929) );
  NAND2XL U19109 ( .A(n19216), .B(w1[37]), .Y(n7927) );
  NAND2XL U19110 ( .A(n3120), .B(y20[5]), .Y(n7926) );
  AOI22XL U19111 ( .A0(n19346), .A1(y10[5]), .B0(n3062), .B1(temp1[5]), .Y(
        n7930) );
  OAI21XL U19112 ( .A0(n19237), .A1(n26588), .B0(n7930), .Y(n8407) );
  NOR2XL U19113 ( .A(n8420), .B(n8407), .Y(n7946) );
  NOR2XL U19114 ( .A(n7931), .B(n7946), .Y(n7943) );
  NAND2XL U19115 ( .A(n6217), .B(y10[6]), .Y(n7935) );
  NAND2XL U19116 ( .A(n19346), .B(w2[6]), .Y(n7934) );
  NAND2XL U19117 ( .A(n3026), .B(w1[38]), .Y(n7933) );
  NAND2XL U19118 ( .A(n3120), .B(y20[6]), .Y(n7932) );
  AOI22XL U19119 ( .A0(n19346), .A1(y10[6]), .B0(n3026), .B1(temp1[6]), .Y(
        n7936) );
  OAI21XL U19120 ( .A0(n19237), .A1(n26587), .B0(n7936), .Y(n8354) );
  NOR2XL U19121 ( .A(n8378), .B(n8354), .Y(n7942) );
  NAND2XL U19122 ( .A(n6217), .B(y10[7]), .Y(n7940) );
  NAND2XL U19123 ( .A(n19346), .B(w2[7]), .Y(n7939) );
  NAND2XL U19124 ( .A(n19161), .B(w1[39]), .Y(n7938) );
  NAND2XL U19125 ( .A(n3120), .B(y20[7]), .Y(n7937) );
  AOI22XL U19126 ( .A0(n19346), .A1(y10[7]), .B0(n3062), .B1(temp1[7]), .Y(
        n7941) );
  OAI21XL U19127 ( .A0(n19237), .A1(n26586), .B0(n7941), .Y(n8356) );
  NOR2XL U19128 ( .A(n8401), .B(n8356), .Y(n7949) );
  NOR2X1 U19129 ( .A(n7942), .B(n7949), .Y(n7952) );
  NAND2XL U19130 ( .A(n7943), .B(n7952), .Y(n7954) );
  NAND2XL U19131 ( .A(n8474), .B(n8427), .Y(n7945) );
  NAND2XL U19132 ( .A(n8420), .B(n8407), .Y(n7944) );
  OAI21XL U19133 ( .A0(n7946), .A1(n7945), .B0(n7944), .Y(n7951) );
  NAND2XL U19134 ( .A(n8378), .B(n8354), .Y(n7948) );
  NAND2XL U19135 ( .A(n8401), .B(n8356), .Y(n7947) );
  OAI21XL U19136 ( .A0(n7949), .A1(n7948), .B0(n7947), .Y(n7950) );
  NAND2XL U19137 ( .A(n6217), .B(y10[8]), .Y(n7959) );
  NAND2XL U19138 ( .A(n19346), .B(w2[8]), .Y(n7958) );
  NAND2XL U19139 ( .A(n19161), .B(w1[40]), .Y(n7957) );
  NAND2XL U19140 ( .A(n3120), .B(y20[8]), .Y(n7956) );
  AOI22XL U19141 ( .A0(n19346), .A1(y10[8]), .B0(n3062), .B1(temp1[8]), .Y(
        n7960) );
  OAI21XL U19142 ( .A0(n19237), .A1(n26585), .B0(n7960), .Y(n8253) );
  NOR2XL U19143 ( .A(n8326), .B(n8253), .Y(n7966) );
  NAND2XL U19144 ( .A(n6217), .B(y10[9]), .Y(n7964) );
  NAND2XL U19145 ( .A(n3027), .B(w2[9]), .Y(n7963) );
  NAND2XL U19146 ( .A(n19161), .B(w1[41]), .Y(n7962) );
  NAND2XL U19147 ( .A(n3120), .B(y20[9]), .Y(n7961) );
  AOI22XL U19148 ( .A0(n19346), .A1(y10[9]), .B0(n3062), .B1(temp1[9]), .Y(
        n7965) );
  OAI21XL U19149 ( .A0(n19237), .A1(n26584), .B0(n7965), .Y(n8255) );
  NOR2XL U19150 ( .A(n8349), .B(n8255), .Y(n8005) );
  NOR2XL U19151 ( .A(n7966), .B(n8005), .Y(n7978) );
  NAND2XL U19152 ( .A(n6217), .B(y10[11]), .Y(n7970) );
  NAND2XL U19153 ( .A(n19346), .B(w2[11]), .Y(n7969) );
  NAND2XL U19154 ( .A(n19161), .B(w1[43]), .Y(n7968) );
  NAND2XL U19155 ( .A(n8104), .B(y20[11]), .Y(n7967) );
  INVX1 U19156 ( .A(n8264), .Y(n8666) );
  AOI22XL U19157 ( .A0(n19346), .A1(y10[11]), .B0(n3026), .B1(temp1[11]), .Y(
        n7971) );
  OAI21XL U19158 ( .A0(n19237), .A1(n26582), .B0(n7971), .Y(n8263) );
  NAND2XL U19159 ( .A(n6217), .B(y10[10]), .Y(n7975) );
  NAND2XL U19160 ( .A(n19346), .B(w2[10]), .Y(n7974) );
  NAND2XL U19161 ( .A(n19161), .B(w1[42]), .Y(n7973) );
  NAND2XL U19162 ( .A(n3120), .B(y20[10]), .Y(n7972) );
  AOI22XL U19163 ( .A0(n3027), .A1(y10[10]), .B0(n19216), .B1(temp1[10]), .Y(
        n7976) );
  OAI21XL U19164 ( .A0(n19237), .A1(n26583), .B0(n7976), .Y(n8260) );
  NOR2XL U19165 ( .A(n8659), .B(n8260), .Y(n7977) );
  NAND2XL U19166 ( .A(n19346), .B(w2[12]), .Y(n7981) );
  NAND2XL U19167 ( .A(n19161), .B(w1[44]), .Y(n7980) );
  NAND2XL U19168 ( .A(n8104), .B(y20[12]), .Y(n7979) );
  AOI22XL U19169 ( .A0(n19346), .A1(y10[12]), .B0(n3026), .B1(temp1[12]), .Y(
        n7983) );
  OAI21XL U19170 ( .A0(n3063), .A1(n26581), .B0(n7983), .Y(n8234) );
  NOR2XL U19171 ( .A(n8674), .B(n8234), .Y(n7989) );
  NAND2XL U19172 ( .A(n6217), .B(y10[13]), .Y(n7987) );
  NAND2XL U19173 ( .A(n3027), .B(w2[13]), .Y(n7986) );
  NAND2XL U19174 ( .A(n19161), .B(w1[45]), .Y(n7985) );
  NAND2XL U19175 ( .A(n8104), .B(y20[13]), .Y(n7984) );
  INVX1 U19176 ( .A(n8237), .Y(n8681) );
  AOI22XL U19177 ( .A0(n19346), .A1(y10[13]), .B0(n3026), .B1(temp1[13]), .Y(
        n7988) );
  OAI21XL U19178 ( .A0(n19237), .A1(n26580), .B0(n7988), .Y(n8236) );
  NAND2XL U19179 ( .A(n6217), .B(y10[15]), .Y(n7993) );
  NAND2XL U19180 ( .A(n19346), .B(w2[15]), .Y(n7992) );
  NAND2XL U19181 ( .A(n3062), .B(w1[47]), .Y(n7991) );
  NAND2XL U19182 ( .A(n8104), .B(y20[15]), .Y(n7990) );
  AOI22XL U19183 ( .A0(n19346), .A1(y10[15]), .B0(n3026), .B1(temp1[15]), .Y(
        n7994) );
  OAI21XL U19184 ( .A0(n19237), .A1(n26578), .B0(n7994), .Y(n8243) );
  NAND2XL U19185 ( .A(n6217), .B(y10[14]), .Y(n7998) );
  NAND2XL U19186 ( .A(n19349), .B(w2[14]), .Y(n7997) );
  NAND2XL U19187 ( .A(n19161), .B(w1[46]), .Y(n7996) );
  NAND2XL U19188 ( .A(n8104), .B(y20[14]), .Y(n7995) );
  INVX1 U19189 ( .A(n8241), .Y(n8686) );
  AOI22XL U19190 ( .A0(n19346), .A1(y10[14]), .B0(n3026), .B1(temp1[14]), .Y(
        n7999) );
  OAI21XL U19191 ( .A0(n19237), .A1(n26579), .B0(n7999), .Y(n8240) );
  NOR2XL U19192 ( .A(n8686), .B(n8240), .Y(n8000) );
  NAND2XL U19193 ( .A(n8326), .B(n8253), .Y(n8004) );
  NAND2XL U19194 ( .A(n8349), .B(n8255), .Y(n8003) );
  NAND2XL U19195 ( .A(n8659), .B(n8260), .Y(n8007) );
  NAND2XL U19196 ( .A(n8666), .B(n8263), .Y(n8006) );
  OAI21XL U19197 ( .A0(n8008), .A1(n8007), .B0(n8006), .Y(n8009) );
  AOI21XL U19198 ( .A0(n8011), .A1(n8010), .B0(n8009), .Y(n8023) );
  NAND2XL U19199 ( .A(n8674), .B(n8234), .Y(n8013) );
  NAND2XL U19200 ( .A(n8681), .B(n8236), .Y(n8012) );
  OAI21XL U19201 ( .A0(n8014), .A1(n8013), .B0(n8012), .Y(n8019) );
  NAND2XL U19202 ( .A(n8686), .B(n8240), .Y(n8016) );
  NAND2XL U19203 ( .A(n8691), .B(n8243), .Y(n8015) );
  OAI21XL U19204 ( .A0(n8017), .A1(n8016), .B0(n8015), .Y(n8018) );
  AOI21XL U19205 ( .A0(n8020), .A1(n8019), .B0(n8018), .Y(n8021) );
  AOI21X1 U19206 ( .A0(n8026), .A1(n8025), .B0(n8024), .Y(n8160) );
  NAND2XL U19207 ( .A(n6217), .B(y10[16]), .Y(n8030) );
  NAND2XL U19208 ( .A(n19349), .B(w2[16]), .Y(n8029) );
  NAND2XL U19209 ( .A(n19161), .B(w1[48]), .Y(n8028) );
  NAND2XL U19210 ( .A(n8104), .B(y20[16]), .Y(n8027) );
  AOI22XL U19211 ( .A0(n19346), .A1(y10[16]), .B0(n3026), .B1(temp1[16]), .Y(
        n8031) );
  OAI21XL U19212 ( .A0(n3063), .A1(n26577), .B0(n8031), .Y(n8306) );
  NOR2XL U19213 ( .A(n8712), .B(n8306), .Y(n8037) );
  NAND2XL U19214 ( .A(n6217), .B(y10[17]), .Y(n8035) );
  NAND2XL U19215 ( .A(n19349), .B(w2[17]), .Y(n8034) );
  NAND2XL U19216 ( .A(n19161), .B(w1[49]), .Y(n8033) );
  NAND2XL U19217 ( .A(n8104), .B(y20[17]), .Y(n8032) );
  AOI22XL U19218 ( .A0(n3027), .A1(y10[17]), .B0(n3026), .B1(temp1[17]), .Y(
        n8036) );
  OAI21XL U19219 ( .A0(n3063), .A1(n26576), .B0(n8036), .Y(n8308) );
  NAND2XL U19220 ( .A(n6217), .B(y10[19]), .Y(n8041) );
  NAND2XL U19221 ( .A(n19349), .B(w2[19]), .Y(n8040) );
  NAND2XL U19222 ( .A(n3026), .B(w1[51]), .Y(n8039) );
  NAND2XL U19223 ( .A(n8104), .B(y20[19]), .Y(n8038) );
  NAND4X1 U19224 ( .A(n8041), .B(n8040), .C(n8039), .D(n8038), .Y(n8316) );
  AOI22XL U19225 ( .A0(n3027), .A1(y10[19]), .B0(n3026), .B1(temp1[19]), .Y(
        n8042) );
  OAI21XL U19226 ( .A0(n3063), .A1(n26574), .B0(n8042), .Y(n8315) );
  NAND2XL U19227 ( .A(n19349), .B(w2[18]), .Y(n8045) );
  NAND2XL U19228 ( .A(n19161), .B(w1[50]), .Y(n8044) );
  NAND2XL U19229 ( .A(n8104), .B(y20[18]), .Y(n8043) );
  AOI22XL U19230 ( .A0(n19346), .A1(y10[18]), .B0(n3026), .B1(temp1[18]), .Y(
        n8047) );
  OAI21XL U19231 ( .A0(n3063), .A1(n26575), .B0(n8047), .Y(n8312) );
  NOR2XL U19232 ( .A(n8788), .B(n8312), .Y(n8048) );
  NAND2XL U19233 ( .A(n6217), .B(y10[20]), .Y(n8053) );
  NAND2XL U19234 ( .A(n19349), .B(w2[20]), .Y(n8052) );
  NAND2XL U19235 ( .A(n3026), .B(w1[52]), .Y(n8051) );
  NAND2XL U19236 ( .A(n8104), .B(y20[20]), .Y(n8050) );
  NAND4X1 U19237 ( .A(n8053), .B(n8052), .C(n8051), .D(n8050), .Y(n8297) );
  INVX1 U19238 ( .A(n8297), .Y(n8798) );
  AOI22XL U19239 ( .A0(n19346), .A1(y10[20]), .B0(n3026), .B1(temp1[20]), .Y(
        n8054) );
  OAI21XL U19240 ( .A0(n3063), .A1(n26573), .B0(n8054), .Y(n8296) );
  NOR2XL U19241 ( .A(n8798), .B(n8296), .Y(n8060) );
  NAND2XL U19242 ( .A(n6217), .B(y10[21]), .Y(n8058) );
  NAND2XL U19243 ( .A(n19349), .B(w2[21]), .Y(n8057) );
  NAND2XL U19244 ( .A(n19216), .B(w1[53]), .Y(n8056) );
  NAND2XL U19245 ( .A(n3120), .B(y20[21]), .Y(n8055) );
  NAND4X1 U19246 ( .A(n8058), .B(n8057), .C(n8056), .D(n8055), .Y(n8299) );
  INVX1 U19247 ( .A(n8299), .Y(n8803) );
  AOI22XL U19248 ( .A0(n3027), .A1(y10[21]), .B0(n3026), .B1(temp1[21]), .Y(
        n8059) );
  OAI21XL U19249 ( .A0(n19237), .A1(n26572), .B0(n8059), .Y(n8298) );
  NAND2XL U19250 ( .A(n6217), .B(y10[23]), .Y(n8064) );
  NAND2XL U19251 ( .A(n19161), .B(w1[55]), .Y(n8062) );
  INVX1 U19252 ( .A(n8196), .Y(n8067) );
  NAND2XL U19253 ( .A(n6217), .B(y10[22]), .Y(n8071) );
  NAND2XL U19254 ( .A(n19349), .B(w2[22]), .Y(n8070) );
  NAND2XL U19255 ( .A(n19161), .B(w1[54]), .Y(n8069) );
  NAND2XL U19256 ( .A(n8104), .B(y20[22]), .Y(n8068) );
  NAND4X1 U19257 ( .A(n8071), .B(n8070), .C(n8069), .D(n8068), .Y(n8303) );
  INVX1 U19258 ( .A(n8303), .Y(n8808) );
  AOI22XL U19259 ( .A0(n3027), .A1(y10[22]), .B0(n3026), .B1(temp1[22]), .Y(
        n8072) );
  OAI21XL U19260 ( .A0(n19237), .A1(n26571), .B0(n8072), .Y(n8302) );
  NOR2XL U19261 ( .A(n8808), .B(n8302), .Y(n8073) );
  NAND2XL U19262 ( .A(n6217), .B(y10[24]), .Y(n8079) );
  NAND2XL U19263 ( .A(n19161), .B(w1[56]), .Y(n8078) );
  AOI22XL U19264 ( .A0(y10[24]), .A1(n19346), .B0(n19161), .B1(temp1[24]), .Y(
        n8080) );
  NAND2XL U19265 ( .A(n6217), .B(y10[25]), .Y(n8084) );
  NAND2XL U19266 ( .A(n3062), .B(w1[57]), .Y(n8082) );
  NAND4X1 U19267 ( .A(n8084), .B(n8083), .C(n8082), .D(n8081), .Y(n8204) );
  INVX1 U19268 ( .A(n8204), .Y(n8171) );
  AOI22XL U19269 ( .A0(y10[25]), .A1(n19346), .B0(n19161), .B1(temp1[25]), .Y(
        n8085) );
  NAND2XL U19270 ( .A(n6217), .B(y10[27]), .Y(n8090) );
  NAND2XL U19271 ( .A(n19161), .B(w1[59]), .Y(n8088) );
  AOI22XL U19272 ( .A0(y10[27]), .A1(n19346), .B0(n19161), .B1(temp1[27]), .Y(
        n8091) );
  NAND2XL U19273 ( .A(n6217), .B(y10[26]), .Y(n8095) );
  NAND2XL U19274 ( .A(n3062), .B(w1[58]), .Y(n8093) );
  INVX1 U19275 ( .A(n8208), .Y(n8169) );
  AOI22XL U19276 ( .A0(y10[26]), .A1(n19346), .B0(n19161), .B1(temp1[26]), .Y(
        n8096) );
  NAND2XL U19277 ( .A(n6217), .B(y10[28]), .Y(n8102) );
  NAND2XL U19278 ( .A(n3062), .B(w1[60]), .Y(n8100) );
  AOI22XL U19279 ( .A0(y10[28]), .A1(n19235), .B0(n19161), .B1(temp1[28]), .Y(
        n8103) );
  NAND2XL U19280 ( .A(n6217), .B(y10[29]), .Y(n8108) );
  NAND2XL U19281 ( .A(n19161), .B(w1[61]), .Y(n8106) );
  OR2X2 U19282 ( .A(n8148), .B(n8192), .Y(n8150) );
  NAND2XL U19283 ( .A(n8712), .B(n8306), .Y(n8115) );
  NAND2XL U19284 ( .A(n8772), .B(n8308), .Y(n8114) );
  OAI21XL U19285 ( .A0(n8116), .A1(n8115), .B0(n8114), .Y(n8121) );
  NAND2XL U19286 ( .A(n8788), .B(n8312), .Y(n8118) );
  NAND2XL U19287 ( .A(n8793), .B(n8315), .Y(n8117) );
  OAI21XL U19288 ( .A0(n8119), .A1(n8118), .B0(n8117), .Y(n8120) );
  AOI21XL U19289 ( .A0(n8122), .A1(n8121), .B0(n8120), .Y(n8134) );
  NAND2XL U19290 ( .A(n8798), .B(n8296), .Y(n8124) );
  NAND2XL U19291 ( .A(n8803), .B(n8298), .Y(n8123) );
  OAI21XL U19292 ( .A0(n8125), .A1(n8124), .B0(n8123), .Y(n8130) );
  NAND2XL U19293 ( .A(n8808), .B(n8302), .Y(n8127) );
  NAND2XL U19294 ( .A(n8067), .B(n8195), .Y(n8126) );
  OAI21XL U19295 ( .A0(n8128), .A1(n8127), .B0(n8126), .Y(n8129) );
  NAND2XL U19296 ( .A(n8135), .B(n8199), .Y(n8137) );
  NAND2XL U19297 ( .A(n8171), .B(n8203), .Y(n8136) );
  OAI21XL U19298 ( .A0(n8138), .A1(n8137), .B0(n8136), .Y(n8143) );
  NAND2XL U19299 ( .A(n8169), .B(n8207), .Y(n8140) );
  NAND2XL U19300 ( .A(n8167), .B(n8180), .Y(n8139) );
  OAI21XL U19301 ( .A0(n8141), .A1(n8140), .B0(n8139), .Y(n8142) );
  AOI21XL U19302 ( .A0(n8144), .A1(n8143), .B0(n8142), .Y(n8154) );
  NAND2XL U19303 ( .A(n8165), .B(n8184), .Y(n8146) );
  NAND2XL U19304 ( .A(n8163), .B(n8188), .Y(n8145) );
  OAI21XL U19305 ( .A0(n8147), .A1(n8146), .B0(n8145), .Y(n8151) );
  INVX8 U19306 ( .A(n3017), .Y(n8482) );
  OAI21X2 U19307 ( .A0(n8482), .A1(n8163), .B0(n8162), .Y(n23844) );
  OAI21X2 U19308 ( .A0(n8482), .A1(n8165), .B0(n8164), .Y(n20374) );
  OAI21X2 U19309 ( .A0(n8482), .A1(n8135), .B0(n8172), .Y(n23870) );
  OAI21X2 U19310 ( .A0(n8482), .A1(n8067), .B0(n8173), .Y(n23760) );
  CMPR22X1 U19311 ( .A(n23844), .B(n8174), .CO(n8992), .S(n23845) );
  CMPR22X1 U19312 ( .A(n20374), .B(n8175), .CO(n8174), .S(n9035) );
  CMPR22X1 U19313 ( .A(n23858), .B(n8176), .CO(n8175), .S(n23859) );
  NAND2XL U19314 ( .A(n3040), .B(n8181), .Y(n8182) );
  INVXL U19315 ( .A(n8188), .Y(n8191) );
  NOR2XL U19316 ( .A(n23185), .B(n23184), .Y(n8212) );
  INVXL U19317 ( .A(n8203), .Y(n8206) );
  NAND2X1 U19318 ( .A(n8482), .B(n8204), .Y(n8205) );
  NAND4X1 U19319 ( .A(n8221), .B(n8220), .C(n8219), .D(n8218), .Y(n23177) );
  INVX1 U19320 ( .A(n23185), .Y(n8233) );
  INVXL U19321 ( .A(n8270), .Y(n8225) );
  INVXL U19322 ( .A(n8228), .Y(n8230) );
  NAND2XL U19323 ( .A(n8230), .B(n8229), .Y(n8232) );
  XNOR2X1 U19324 ( .A(n23760), .B(n8233), .Y(n8259) );
  NAND2XL U19325 ( .A(n3092), .B(n8238), .Y(n8239) );
  OAI21XL U19326 ( .A0(n3092), .A1(n8590), .B0(n8239), .Y(n8351) );
  INVXL U19327 ( .A(n8240), .Y(n8687) );
  OAI21XL U19328 ( .A0(n3040), .A1(n8687), .B0(n8242), .Y(n8569) );
  INVXL U19329 ( .A(n8243), .Y(n8692) );
  OAI21XL U19330 ( .A0(n3040), .A1(n8692), .B0(n8245), .Y(n8560) );
  NAND2XL U19331 ( .A(n3092), .B(n8560), .Y(n8246) );
  OAI21XL U19332 ( .A0(n3092), .A1(n8247), .B0(n8246), .Y(n8370) );
  INVXL U19333 ( .A(n8370), .Y(n8248) );
  NAND2XL U19334 ( .A(n3162), .B(n8248), .Y(n8249) );
  OAI21XL U19335 ( .A0(n3162), .A1(n8351), .B0(n8249), .Y(n8462) );
  INVXL U19336 ( .A(n8267), .Y(n8250) );
  NAND2XL U19337 ( .A(n8250), .B(n8269), .Y(n8251) );
  XOR2X1 U19338 ( .A(n8252), .B(n8251), .Y(n8405) );
  OAI21XL U19339 ( .A0(n3040), .A1(n8350), .B0(n8257), .Y(n8576) );
  NAND2XL U19340 ( .A(n3092), .B(n8576), .Y(n8258) );
  OAI21XL U19341 ( .A0(n3092), .A1(n8536), .B0(n8258), .Y(n8359) );
  INVXL U19342 ( .A(n8260), .Y(n8660) );
  OAI21XL U19343 ( .A0(n3040), .A1(n8660), .B0(n8262), .Y(n8531) );
  INVXL U19344 ( .A(n8263), .Y(n8667) );
  OAI21XL U19345 ( .A0(n3040), .A1(n8667), .B0(n8265), .Y(n8559) );
  AOI22XL U19346 ( .A0(n8592), .A1(n8531), .B0(n3092), .B1(n8559), .Y(n8353)
         );
  NAND2XL U19347 ( .A(n3162), .B(n8353), .Y(n8266) );
  OAI21XL U19348 ( .A0(n3162), .A1(n8359), .B0(n8266), .Y(n8467) );
  OAI22XL U19349 ( .A0(n8462), .A1(n8434), .B0(n3157), .B1(n8467), .Y(n8489)
         );
  NOR2XL U19350 ( .A(n8267), .B(n8270), .Y(n8273) );
  OAI21XL U19351 ( .A0(n8270), .A1(n8269), .B0(n8268), .Y(n8271) );
  OAI21XL U19352 ( .A0(n8294), .A1(n8290), .B0(n8291), .Y(n8278) );
  NAND2X2 U19353 ( .A(n8565), .B(n8289), .Y(n8614) );
  INVXL U19354 ( .A(n8290), .Y(n8292) );
  OAI21XL U19355 ( .A0(n3040), .A1(n8804), .B0(n8300), .Y(n8554) );
  NAND2XL U19356 ( .A(n3092), .B(n8554), .Y(n8301) );
  INVXL U19357 ( .A(n8302), .Y(n8809) );
  OAI21XL U19358 ( .A0(n3040), .A1(n8809), .B0(n8304), .Y(n8553) );
  NAND2XL U19359 ( .A(n3162), .B(n8372), .Y(n8305) );
  OAI21XL U19360 ( .A0(n8606), .A1(n8363), .B0(n8305), .Y(n8669) );
  INVXL U19361 ( .A(n8669), .Y(n8322) );
  CLKINVX3 U19362 ( .A(n8405), .Y(n8434) );
  OAI21XL U19363 ( .A0(n3040), .A1(n8773), .B0(n8310), .Y(n8524) );
  NAND2XL U19364 ( .A(n3092), .B(n8524), .Y(n8311) );
  OAI21XL U19365 ( .A0(n3092), .A1(n8586), .B0(n8311), .Y(n8367) );
  OAI21XL U19366 ( .A0(n3040), .A1(n8789), .B0(n8314), .Y(n8552) );
  NAND2XL U19367 ( .A(n3092), .B(n8534), .Y(n8318) );
  OAI21XL U19368 ( .A0(n3092), .A1(n8319), .B0(n8318), .Y(n8366) );
  INVXL U19369 ( .A(n8366), .Y(n8320) );
  NAND2XL U19370 ( .A(n3162), .B(n8320), .Y(n8321) );
  OAI21XL U19371 ( .A0(n3162), .A1(n8367), .B0(n8321), .Y(n8463) );
  AOI22XL U19372 ( .A0(n8592), .A1(n8576), .B0(n3092), .B1(n8531), .Y(n8394)
         );
  NAND2XL U19373 ( .A(n3092), .B(n8328), .Y(n8329) );
  OAI21XL U19374 ( .A0(n3092), .A1(n8330), .B0(n8329), .Y(n8390) );
  INVXL U19375 ( .A(n8390), .Y(n8331) );
  AOI22XL U19376 ( .A0(n4591), .A1(n8394), .B0(n8331), .B1(n8606), .Y(n8412)
         );
  NAND2XL U19377 ( .A(n3092), .B(n8569), .Y(n8332) );
  OAI21XL U19378 ( .A0(n3092), .A1(n8557), .B0(n8332), .Y(n8387) );
  AOI22XL U19379 ( .A0(n8592), .A1(n8560), .B0(n3092), .B1(n8333), .Y(n8382)
         );
  NAND2XL U19380 ( .A(n3162), .B(n8382), .Y(n8334) );
  OAI21XL U19381 ( .A0(n3162), .A1(n8387), .B0(n8334), .Y(n8404) );
  NAND2XL U19382 ( .A(n3092), .B(n8553), .Y(n8335) );
  OAI21XL U19383 ( .A0(n3092), .A1(n8336), .B0(n8335), .Y(n8383) );
  OAI21XL U19384 ( .A0(n8606), .A1(n8383), .B0(n8337), .Y(n8676) );
  INVXL U19385 ( .A(n8676), .Y(n8345) );
  NAND2XL U19386 ( .A(n3092), .B(n8552), .Y(n8338) );
  OAI21XL U19387 ( .A0(n3092), .A1(n8339), .B0(n8338), .Y(n8380) );
  NAND2XL U19388 ( .A(n3092), .B(n8340), .Y(n8341) );
  OAI21XL U19389 ( .A0(n8259), .A1(n8342), .B0(n8341), .Y(n8386) );
  INVXL U19390 ( .A(n8386), .Y(n8343) );
  NAND2XL U19391 ( .A(n3162), .B(n8343), .Y(n8344) );
  AOI22XL U19392 ( .A0(n8502), .A1(n3086), .B0(n8503), .B1(n3154), .Y(n8346)
         );
  INVXL U19393 ( .A(n8351), .Y(n8352) );
  AOI22XL U19394 ( .A0(n4591), .A1(n8353), .B0(n8352), .B1(n8606), .Y(n8435)
         );
  OAI21XL U19395 ( .A0(n8482), .A1(n8402), .B0(n8358), .Y(n8540) );
  AOI22XL U19396 ( .A0(n8592), .A1(n8573), .B0(n3092), .B1(n8540), .Y(n8464)
         );
  INVXL U19397 ( .A(n8464), .Y(n8362) );
  INVXL U19398 ( .A(n8359), .Y(n8360) );
  NAND2XL U19399 ( .A(n3162), .B(n8360), .Y(n8361) );
  OAI21XL U19400 ( .A0(n3162), .A1(n8362), .B0(n8361), .Y(n8431) );
  INVXL U19401 ( .A(n8363), .Y(n8364) );
  NAND2XL U19402 ( .A(n3162), .B(n8364), .Y(n8365) );
  OAI21XL U19403 ( .A0(n3162), .A1(n8366), .B0(n8365), .Y(n8436) );
  INVXL U19404 ( .A(n8436), .Y(n8371) );
  INVXL U19405 ( .A(n8367), .Y(n8368) );
  NAND2XL U19406 ( .A(n3162), .B(n8368), .Y(n8369) );
  OAI21XL U19407 ( .A0(n3162), .A1(n8370), .B0(n8369), .Y(n8433) );
  NAND2XL U19408 ( .A(n8434), .B(n4591), .Y(n8555) );
  INVXL U19409 ( .A(n8380), .Y(n8381) );
  AOI22XL U19410 ( .A0(n8447), .A1(n8382), .B0(n8381), .B1(n8606), .Y(n8452)
         );
  INVXL U19411 ( .A(n8383), .Y(n8384) );
  NAND2XL U19412 ( .A(n3162), .B(n8384), .Y(n8385) );
  OAI21XL U19413 ( .A0(n3162), .A1(n8386), .B0(n8385), .Y(n8453) );
  INVXL U19414 ( .A(n8387), .Y(n8388) );
  NAND2XL U19415 ( .A(n3162), .B(n8388), .Y(n8389) );
  OAI21XL U19416 ( .A0(n3162), .A1(n8390), .B0(n8389), .Y(n8451) );
  NAND2XL U19417 ( .A(n3092), .B(n8391), .Y(n8392) );
  OAI21XL U19418 ( .A0(n3092), .A1(n8393), .B0(n8392), .Y(n8410) );
  NAND2XL U19419 ( .A(n3162), .B(n8394), .Y(n8395) );
  OAI21XL U19420 ( .A0(n3162), .A1(n8410), .B0(n8395), .Y(n8448) );
  CLKINVX2 U19421 ( .A(n8610), .Y(n8593) );
  OAI21XL U19422 ( .A0(n8613), .A1(n3154), .B0(n8593), .Y(n8396) );
  OAI22XL U19423 ( .A0(n8406), .A1(n3087), .B0(n8405), .B1(n8404), .Y(n8678)
         );
  INVX1 U19424 ( .A(n8606), .Y(n8447) );
  OAI21XL U19425 ( .A0(n8482), .A1(n8421), .B0(n8409), .Y(n8564) );
  AOI22XL U19426 ( .A0(n8592), .A1(n8564), .B0(n3092), .B1(n8573), .Y(n8446)
         );
  INVXL U19427 ( .A(n8410), .Y(n8411) );
  AOI22XL U19428 ( .A0(n8447), .A1(n8446), .B0(n8411), .B1(n8606), .Y(n8499)
         );
  OAI21XL U19429 ( .A0(n8678), .A1(n3086), .B0(n8414), .Y(n8415) );
  OAI21XL U19430 ( .A0(n8482), .A1(n8460), .B0(n8426), .Y(n8544) );
  AOI22XL U19431 ( .A0(n8592), .A1(n8562), .B0(n3092), .B1(n8544), .Y(n8483)
         );
  NAND2XL U19432 ( .A(n3092), .B(n8564), .Y(n8429) );
  OAI21XL U19433 ( .A0(n3092), .A1(n8542), .B0(n8429), .Y(n8466) );
  INVXL U19434 ( .A(n8466), .Y(n8430) );
  AOI22XL U19435 ( .A0(n8447), .A1(n8483), .B0(n8430), .B1(n8606), .Y(n8514)
         );
  AOI21XL U19436 ( .A0(n8432), .A1(n8601), .B0(n8610), .Y(n8439) );
  NAND2XL U19437 ( .A(n8655), .B(n3154), .Y(n8438) );
  AOI2BB2X1 U19438 ( .B0(n8437), .B1(n3157), .A0N(n3157), .A1N(n8436), .Y(
        n8654) );
  OAI21XL U19439 ( .A0(n3160), .A1(n8442), .B0(n8441), .Y(n8627) );
  NOR2XL U19440 ( .A(n8627), .B(n8626), .Y(n8897) );
  INVXL U19441 ( .A(n8897), .Y(n8902) );
  INVXL U19442 ( .A(n8542), .Y(n8445) );
  AOI22XL U19443 ( .A0(n8592), .A1(n8544), .B0(n3092), .B1(n8445), .Y(n8498)
         );
  AOI22XL U19444 ( .A0(n8447), .A1(n8498), .B0(n8446), .B1(n8606), .Y(n8608)
         );
  INVXL U19445 ( .A(n8448), .Y(n8449) );
  AOI22XL U19446 ( .A0(n8608), .A1(n3087), .B0(n8449), .B1(n3157), .Y(n8450)
         );
  AOI21XL U19447 ( .A0(n8450), .A1(n8601), .B0(n8610), .Y(n8455) );
  NAND2XL U19448 ( .A(n8662), .B(n3154), .Y(n8454) );
  NAND2XL U19449 ( .A(n4591), .B(n8592), .Y(n8571) );
  INVXL U19450 ( .A(n8571), .Y(n8550) );
  AOI22XL U19451 ( .A0(n8455), .A1(n8454), .B0(n8790), .B1(n8610), .Y(n8456)
         );
  AOI21XL U19452 ( .A0(n8458), .A1(n8823), .B0(n3155), .Y(n8457) );
  OAI21XL U19453 ( .A0(n3160), .A1(n8458), .B0(n8457), .Y(n8629) );
  NAND2XL U19454 ( .A(n8902), .B(n8461), .Y(n8891) );
  OAI22XL U19455 ( .A0(n8463), .A1(n3087), .B0(n3157), .B1(n8462), .Y(n8671)
         );
  NAND2XL U19456 ( .A(n3162), .B(n8464), .Y(n8465) );
  OAI21XL U19457 ( .A0(n3162), .A1(n8466), .B0(n8465), .Y(n8484) );
  OAI22XL U19458 ( .A0(n8671), .A1(n3086), .B0(n8468), .B1(n3154), .Y(n8469)
         );
  NAND2XL U19459 ( .A(n8469), .B(n8593), .Y(n8470) );
  OAI21XL U19460 ( .A0(n8795), .A1(n8593), .B0(n8470), .Y(n8471) );
  AOI21XL U19461 ( .A0(n8473), .A1(n8823), .B0(n3155), .Y(n8472) );
  OAI21XL U19462 ( .A0(n3160), .A1(n8473), .B0(n8472), .Y(n8633) );
  NOR2XL U19463 ( .A(n8633), .B(n8632), .Y(n8892) );
  NOR2XL U19464 ( .A(n8891), .B(n8892), .Y(n8635) );
  INVXL U19465 ( .A(n8709), .Y(n8491) );
  OAI21XL U19466 ( .A0(n8482), .A1(n8510), .B0(n8481), .Y(n8579) );
  AOI22XL U19467 ( .A0(n8592), .A1(n8578), .B0(n8259), .B1(n8579), .Y(n8513)
         );
  AOI22XL U19468 ( .A0(n4591), .A1(n8513), .B0(n8483), .B1(n8606), .Y(n8486)
         );
  INVXL U19469 ( .A(n8484), .Y(n8485) );
  AOI22XL U19470 ( .A0(n8486), .A1(n8434), .B0(n8485), .B1(n3157), .Y(n8487)
         );
  AOI21XL U19471 ( .A0(n8487), .A1(n8601), .B0(n8610), .Y(n8488) );
  OAI21XL U19472 ( .A0(n3086), .A1(n8489), .B0(n8488), .Y(n8490) );
  OAI21XL U19473 ( .A0(n8491), .A1(n8593), .B0(n8490), .Y(n8492) );
  NAND2XL U19474 ( .A(n8493), .B(n8492), .Y(n8495) );
  AOI21XL U19475 ( .A0(n8495), .A1(n8823), .B0(n3155), .Y(n8494) );
  OAI21XL U19476 ( .A0(n3160), .A1(n8495), .B0(n8494), .Y(n8620) );
  OR2X2 U19477 ( .A(n8620), .B(n8619), .Y(n8939) );
  AOI22XL U19478 ( .A0(n4591), .A1(n8607), .B0(n8498), .B1(n8606), .Y(n8500)
         );
  AOI22XL U19479 ( .A0(n8500), .A1(n8434), .B0(n8499), .B1(n3157), .Y(n8501)
         );
  AOI21XL U19480 ( .A0(n8501), .A1(n8601), .B0(n8610), .Y(n8505) );
  NAND2XL U19481 ( .A(n8502), .B(n3154), .Y(n8504) );
  AOI22XL U19482 ( .A0(n8505), .A1(n8504), .B0(n8769), .B1(n8610), .Y(n8506)
         );
  AOI21XL U19483 ( .A0(n8508), .A1(n8823), .B0(n3155), .Y(n8507) );
  OAI21XL U19484 ( .A0(n3160), .A1(n8508), .B0(n8507), .Y(n8622) );
  NAND2XL U19485 ( .A(n8939), .B(n8908), .Y(n8625) );
  AOI22XL U19486 ( .A0(n8512), .A1(n3086), .B0(n3154), .B1(n8511), .Y(n8683)
         );
  AOI22XL U19487 ( .A0(n8515), .A1(n3087), .B0(n8514), .B1(n3157), .Y(n8516)
         );
  AOI21XL U19488 ( .A0(n8516), .A1(n3086), .B0(n8610), .Y(n8519) );
  NAND2XL U19489 ( .A(n8517), .B(n3154), .Y(n8518) );
  AOI22XL U19490 ( .A0(n8610), .A1(n8683), .B0(n8519), .B1(n8518), .Y(n8520)
         );
  NOR2XL U19491 ( .A(n8520), .B(n8614), .Y(n8522) );
  NAND2XL U19492 ( .A(n8522), .B(n8668), .Y(n8521) );
  OAI211XL U19493 ( .A0(n9027), .A1(n8522), .B0(n6169), .C0(n8521), .Y(n8523)
         );
  OAI21XL U19494 ( .A0(n3086), .A1(n8551), .B0(n8593), .Y(n8530) );
  NAND2XL U19495 ( .A(n8570), .B(n8524), .Y(n8527) );
  AOI31XL U19496 ( .A0(n8527), .A1(n8526), .A2(n8525), .B0(n8593), .Y(n8529)
         );
  AOI211XL U19497 ( .A0(n8531), .A1(n8530), .B0(n8529), .C0(n8528), .Y(n8549)
         );
  AOI21XL U19498 ( .A0(n3086), .A1(n8592), .B0(n8532), .Y(n8535) );
  INVXL U19499 ( .A(n8570), .Y(n8588) );
  AOI211XL U19500 ( .A0(n3086), .A1(n4591), .B0(n8588), .C0(n8593), .Y(n8533)
         );
  OAI21XL U19501 ( .A0(n8535), .A1(n8534), .B0(n8533), .Y(n8548) );
  NOR2XL U19502 ( .A(n8610), .B(n8537), .Y(n8561) );
  AOI21XL U19503 ( .A0(n8538), .A1(n8447), .B0(n8561), .Y(n8539) );
  OAI21XL U19504 ( .A0(n8541), .A1(n8540), .B0(n8539), .Y(n8547) );
  AOI21XL U19505 ( .A0(n8561), .A1(n8592), .B0(n8542), .Y(n8545) );
  OAI21XL U19506 ( .A0(n3087), .A1(n8447), .B0(n8561), .Y(n8543) );
  OAI21XL U19507 ( .A0(n8545), .A1(n8544), .B0(n8543), .Y(n8546) );
  NAND4XL U19508 ( .A(n8549), .B(n8548), .C(n8547), .D(n8546), .Y(n8600) );
  AOI21XL U19509 ( .A0(n8550), .A1(n8434), .B0(n8601), .Y(n8574) );
  NAND2XL U19510 ( .A(n8601), .B(n8551), .Y(n8563) );
  AOI22XL U19511 ( .A0(n8574), .A1(n8553), .B0(n8563), .B1(n8552), .Y(n8558)
         );
  OAI21XL U19512 ( .A0(n8555), .A1(n8554), .B0(n3154), .Y(n8556) );
  AOI31XL U19513 ( .A0(n8558), .A1(n8557), .A2(n8556), .B0(n8593), .Y(n8568)
         );
  AOI21XL U19514 ( .A0(n8588), .A1(n8447), .B0(n8593), .Y(n8585) );
  NAND2XL U19515 ( .A(n3154), .B(n3157), .Y(n8575) );
  OAI21XL U19516 ( .A0(n8575), .A1(n8447), .B0(n8593), .Y(n8589) );
  AOI22XL U19517 ( .A0(n8585), .A1(n8560), .B0(n8589), .B1(n8559), .Y(n8567)
         );
  INVXL U19518 ( .A(n8561), .Y(n8580) );
  AOI22XL U19519 ( .A0(n8580), .A1(n8564), .B0(n8563), .B1(n8562), .Y(n8566)
         );
  NAND4BXL U19520 ( .AN(n8568), .B(n8567), .C(n8566), .D(n8565), .Y(n8597) );
  OAI211XL U19521 ( .A0(n8571), .A1(n8570), .B0(n8610), .C0(n8569), .Y(n8584)
         );
  AOI22XL U19522 ( .A0(n8574), .A1(n8573), .B0(n8604), .B1(n8606), .Y(n8583)
         );
  INVXL U19523 ( .A(n8575), .Y(n8577) );
  OAI21XL U19524 ( .A0(n8577), .A1(n8610), .B0(n8576), .Y(n8582) );
  OAI22XL U19525 ( .A0(n8580), .A1(n3157), .B0(n8579), .B1(n8578), .Y(n8581)
         );
  NAND4XL U19526 ( .A(n8584), .B(n8583), .C(n8582), .D(n8581), .Y(n8596) );
  INVXL U19527 ( .A(n8585), .Y(n8587) );
  AOI211XL U19528 ( .A0(n8588), .A1(n8592), .B0(n8587), .C0(n8586), .Y(n8595)
         );
  INVXL U19529 ( .A(n8589), .Y(n8591) );
  AOI211XL U19530 ( .A0(n8593), .A1(n8592), .B0(n8591), .C0(n8590), .Y(n8594)
         );
  OR4X2 U19531 ( .A(n8597), .B(n8596), .C(n8595), .D(n8594), .Y(n8599) );
  AOI22XL U19532 ( .A0(n8603), .A1(n3154), .B0(n8602), .B1(n8601), .Y(n8688)
         );
  NAND2XL U19533 ( .A(n8688), .B(n8610), .Y(n8616) );
  INVXL U19534 ( .A(n8604), .Y(n8605) );
  AOI22XL U19535 ( .A0(n3087), .A1(n8609), .B0(n8608), .B1(n3157), .Y(n8611)
         );
  AOI21XL U19536 ( .A0(n8611), .A1(n3086), .B0(n8610), .Y(n8612) );
  OAI21XL U19537 ( .A0(n3086), .A1(n8613), .B0(n8612), .Y(n8615) );
  AOI21XL U19538 ( .A0(n8616), .A1(n8615), .B0(n8614), .Y(n8618) );
  NAND2XL U19539 ( .A(n8618), .B(n8668), .Y(n8617) );
  OAI211XL U19540 ( .A0(n8618), .A1(n9027), .B0(n6169), .C0(n8617), .Y(n8942)
         );
  NAND2XL U19541 ( .A(n8943), .B(n8942), .Y(n8905) );
  NAND2XL U19542 ( .A(n8620), .B(n8619), .Y(n8938) );
  INVXL U19543 ( .A(n8938), .Y(n8906) );
  NAND2XL U19544 ( .A(n8622), .B(n8621), .Y(n8907) );
  INVXL U19545 ( .A(n8907), .Y(n8623) );
  AOI21XL U19546 ( .A0(n8908), .A1(n8906), .B0(n8623), .Y(n8624) );
  INVXL U19547 ( .A(n8901), .Y(n8631) );
  NAND2XL U19548 ( .A(n8629), .B(n8628), .Y(n8898) );
  INVXL U19549 ( .A(n8898), .Y(n8630) );
  OAI21XL U19550 ( .A0(n8890), .A1(n8892), .B0(n8893), .Y(n8634) );
  OAI21XL U19551 ( .A0(n8763), .A1(n8920), .B0(n8764), .Y(n8650) );
  OAI21XL U19552 ( .A0(n3160), .A1(n8665), .B0(n8664), .Y(n8696) );
  OAI21XL U19553 ( .A0(n3157), .A1(n8669), .B0(n3154), .Y(n8670) );
  OAI21XL U19554 ( .A0(n3160), .A1(n8673), .B0(n8672), .Y(n8698) );
  OAI21XL U19555 ( .A0(n3157), .A1(n8676), .B0(n3154), .Y(n8677) );
  OAI21XL U19556 ( .A0(n3160), .A1(n8680), .B0(n8679), .Y(n8700) );
  OAI21XL U19557 ( .A0(n3160), .A1(n8685), .B0(n8684), .Y(n8704) );
  OAI21XL U19558 ( .A0(n3160), .A1(n8690), .B0(n8689), .Y(n8706) );
  OAI21XL U19559 ( .A0(n8749), .A1(n8755), .B0(n8750), .Y(n8742) );
  OAI21XL U19560 ( .A0(n8736), .A1(n8745), .B0(n8737), .Y(n8701) );
  OAI21XL U19561 ( .A0(n8723), .A1(n8728), .B0(n8724), .Y(n8854) );
  AOI21XL U19562 ( .A0(n8860), .A1(n8851), .B0(n8854), .Y(n8707) );
  OAI21XL U19563 ( .A0(n8863), .A1(n8708), .B0(n8707), .Y(n8718) );
  OAI21XL U19564 ( .A0(n3160), .A1(n8711), .B0(n8710), .Y(n8715) );
  OAI21XL U19565 ( .A0(n8863), .A1(n8722), .B0(n8721), .Y(n8727) );
  OAI21XL U19566 ( .A0(n8863), .A1(n8774), .B0(n8781), .Y(n8731) );
  AOI21XL U19567 ( .A0(n8742), .A1(n8746), .B0(n8733), .Y(n8734) );
  OAI21XL U19568 ( .A0(n8863), .A1(n8735), .B0(n8734), .Y(n8740) );
  OAI21XL U19569 ( .A0(n8863), .A1(n8744), .B0(n8743), .Y(n8748) );
  OAI21XL U19570 ( .A0(n8863), .A1(n8754), .B0(n8755), .Y(n8753) );
  OAI21XL U19571 ( .A0(n8760), .A1(n8919), .B0(n8920), .Y(n8761) );
  OAI21XL U19572 ( .A0(n8864), .A1(n8855), .B0(n8865), .Y(n8777) );
  OR2X2 U19573 ( .A(n8870), .B(n8830), .Y(n8834) );
  OAI21XL U19574 ( .A0(n8883), .A1(n8876), .B0(n8884), .Y(n8818) );
  OAI21XL U19575 ( .A0(n8869), .A1(n8830), .B0(n8826), .Y(n8827) );
  OAI21XL U19576 ( .A0(n8882), .A1(n8838), .B0(n8837), .Y(n8841) );
  OAI21XL U19577 ( .A0(n8882), .A1(n8847), .B0(n8848), .Y(n8846) );
  OAI21XL U19578 ( .A0(n8857), .A1(n8856), .B0(n8855), .Y(n8858) );
  OAI21XL U19579 ( .A0(n8863), .A1(n8862), .B0(n8861), .Y(n8868) );
  OAI21XL U19580 ( .A0(n8882), .A1(n8870), .B0(n8869), .Y(n8874) );
  AOI21XL U19581 ( .A0(n8879), .A1(n8878), .B0(n8877), .Y(n8880) );
  OAI21XL U19582 ( .A0(n8882), .A1(n8881), .B0(n8880), .Y(n8887) );
  CMPR22X1 U19583 ( .A(n23816), .B(n8888), .CO(n8176), .S(n23817) );
  INVXL U19584 ( .A(n8889), .Y(n8904) );
  OAI21XL U19585 ( .A0(n8904), .A1(n8897), .B0(n8901), .Y(n8900) );
  XNOR2X1 U19586 ( .A(n8900), .B(n8899), .Y(n20440) );
  XOR2X1 U19587 ( .A(n8904), .B(n8903), .Y(n20443) );
  AOI21XL U19588 ( .A0(n8941), .A1(n8939), .B0(n8906), .Y(n8910) );
  NAND2XL U19589 ( .A(n8908), .B(n8907), .Y(n8909) );
  AOI21XL U19590 ( .A0(n8930), .A1(n8915), .B0(n8911), .Y(n8914) );
  AOI21XL U19591 ( .A0(n8930), .A1(n8918), .B0(n8917), .Y(n8923) );
  OAI21XL U19592 ( .A0(n8927), .A1(n8926), .B0(n8925), .Y(n8928) );
  AOI21XL U19593 ( .A0(n8930), .A1(n8929), .B0(n8928), .Y(n8933) );
  OR2X2 U19594 ( .A(n20411), .B(n20432), .Y(n8969) );
  CMPR22X1 U19595 ( .A(n23810), .B(n8937), .CO(n8888), .S(n23811) );
  NAND2XL U19596 ( .A(n8939), .B(n8938), .Y(n8940) );
  INVXL U19597 ( .A(n8942), .Y(n8944) );
  XNOR2XL U19598 ( .A(n8944), .B(n8943), .Y(n9028) );
  OAI21XL U19599 ( .A0(n8947), .A1(n8946), .B0(n8945), .Y(n8949) );
  AOI31X4 U19600 ( .A0(n8973), .A1(n8952), .A2(n8976), .B0(n8951), .Y(n20473)
         );
  AOI2BB1XL U19601 ( .A0N(n8956), .A1N(n20432), .B0(n20411), .Y(n8957) );
  AOI2BB1XL U19602 ( .A0N(n8957), .A1N(n20461), .B0(n20415), .Y(n8958) );
  AOI2BB1X1 U19603 ( .A0N(n8958), .A1N(n20458), .B0(n20457), .Y(n8959) );
  AOI2BB1X2 U19604 ( .A0N(n8959), .A1N(n20454), .B0(n20453), .Y(n8960) );
  AOI2BB1X2 U19605 ( .A0N(n8960), .A1N(n20450), .B0(n20449), .Y(n8961) );
  AOI2BB1X2 U19606 ( .A0N(n8961), .A1N(n20543), .B0(n20542), .Y(n8962) );
  AOI2BB1X2 U19607 ( .A0N(n8962), .A1N(n20562), .B0(n20561), .Y(n8963) );
  AOI2BB1X2 U19608 ( .A0N(n8963), .A1N(n20400), .B0(n20404), .Y(n8964) );
  AOI2BB1X2 U19609 ( .A0N(n8964), .A1N(n20402), .B0(n9030), .Y(n9009) );
  NAND2XL U19610 ( .A(n23760), .B(n9009), .Y(n8988) );
  OAI21XL U19611 ( .A0(n9016), .A1(n9028), .B0(n8965), .Y(n8966) );
  OAI21XL U19612 ( .A0(n8970), .A1(n8969), .B0(n8968), .Y(n8971) );
  CMPR22X1 U19613 ( .A(n23870), .B(n23760), .CO(n8937), .S(n23872) );
  XOR2X1 U19614 ( .A(n23845), .B(n8982), .Y(n23843) );
  INVXL U19615 ( .A(n9035), .Y(n8983) );
  ADDFHX1 U19616 ( .A(n8988), .B(n3071), .CI(n23872), .CO(n8987), .S(n23869)
         );
  OR4X2 U19617 ( .A(n23815), .B(n23809), .C(n23759), .D(n23869), .Y(n8989) );
  OR4X2 U19618 ( .A(n23843), .B(n9029), .C(n23857), .D(n8989), .Y(n8990) );
  NOR2X1 U19619 ( .A(n23689), .B(n8990), .Y(n8996) );
  CMPR22X1 U19620 ( .A(n23690), .B(n8992), .CO(n8993), .S(n23691) );
  NOR2BX1 U19621 ( .AN(n8994), .B(n8993), .Y(n8995) );
  INVXL U19622 ( .A(n20477), .Y(n9012) );
  NAND4XL U19623 ( .A(n20439), .B(n9016), .C(n9015), .D(n20443), .Y(n9017) );
  INVXL U19624 ( .A(n20440), .Y(n20390) );
  NAND4BXL U19625 ( .AN(n9025), .B(n9024), .C(n20400), .D(n20561), .Y(n9026)
         );
  INVXL U19626 ( .A(n20379), .Y(n9033) );
  AOI22XL U19627 ( .A0(n23873), .A1(n9035), .B0(n23871), .B1(n20374), .Y(n9036) );
  INVXL U19628 ( .A(n24451), .Y(n9039) );
  AND2X1 U19629 ( .A(n23970), .B(n25886), .Y(n25664) );
  INVX1 U19630 ( .A(n8104), .Y(n20748) );
  AOI21XL U19631 ( .A0(n24447), .A1(n24525), .B0(n9040), .Y(n9041) );
  INVXL U19632 ( .A(n9041), .Y(n25859) );
  INVX8 U19633 ( .A(n3223), .Y(n25243) );
  NAND2X4 U19634 ( .A(n4582), .B(n3024), .Y(n22472) );
  INVX4 U19635 ( .A(n22472), .Y(n14417) );
  AOI21XL U19636 ( .A0(n14417), .A1(y11[20]), .B0(n25157), .Y(n9042) );
  NAND2X4 U19637 ( .A(n4580), .B(n6174), .Y(n9053) );
  INVXL U19638 ( .A(n25152), .Y(n9044) );
  INVX8 U19639 ( .A(n9053), .Y(n14427) );
  AOI22XL U19640 ( .A0(n11536), .A1(data[10]), .B0(in_valid_d), .B1(w1[266]), 
        .Y(n9048) );
  NAND2X1 U19641 ( .A(n4826), .B(target_temp[10]), .Y(n11520) );
  OAI211X2 U19642 ( .A0(n23992), .A1(n25243), .B0(n9048), .C0(n11520), .Y(
        M2_b_10_) );
  INVXL U19643 ( .A(n25140), .Y(n9051) );
  AOI2BB2X1 U19644 ( .B0(n9164), .B1(y12[3]), .A0N(n9053), .A1N(n25894), .Y(
        n9055) );
  INVXL U19645 ( .A(n25141), .Y(n9054) );
  AOI22X1 U19646 ( .A0(n25229), .A1(y12[1]), .B0(n14427), .B1(y10[1]), .Y(
        n9057) );
  INVXL U19647 ( .A(n25139), .Y(n9056) );
  AOI22XL U19648 ( .A0(n11536), .A1(data[22]), .B0(in_valid_d), .B1(w1[278]), 
        .Y(n9059) );
  AOI22XL U19649 ( .A0(n9164), .A1(y12[4]), .B0(n14427), .B1(y10[4]), .Y(n9061) );
  INVXL U19650 ( .A(n25142), .Y(n9060) );
  INVXL U19651 ( .A(n25144), .Y(n9065) );
  INVXL U19652 ( .A(learning_rate[18]), .Y(n23988) );
  AOI22XL U19653 ( .A0(n4566), .A1(data[19]), .B0(in_valid_d), .B1(w1[275]), 
        .Y(n9068) );
  INVXL U19654 ( .A(n4771), .Y(n9069) );
  NAND2X1 U19655 ( .A(n14427), .B(y10[17]), .Y(n9072) );
  AOI22XL U19656 ( .A0(n11536), .A1(data[6]), .B0(in_valid_d), .B1(w1[262]), 
        .Y(n9073) );
  NAND2X1 U19657 ( .A(n9164), .B(target_temp[6]), .Y(n11511) );
  INVX1 U19658 ( .A(learning_rate[7]), .Y(n23995) );
  AOI22XL U19659 ( .A0(n11536), .A1(data[7]), .B0(in_valid_d), .B1(w1[263]), 
        .Y(n9074) );
  OAI211X1 U19660 ( .A0(n23995), .A1(n25243), .B0(n9074), .C0(n11504), .Y(
        M2_b_7_) );
  AOI22XL U19661 ( .A0(n25229), .A1(y12[16]), .B0(n14427), .B1(y10[16]), .Y(
        n9076) );
  INVXL U19662 ( .A(n25154), .Y(n9075) );
  AOI22XL U19663 ( .A0(n11536), .A1(data[8]), .B0(in_valid_d), .B1(w1[264]), 
        .Y(n9077) );
  NAND2X1 U19664 ( .A(n4826), .B(target_temp[8]), .Y(n11505) );
  INVXL U19665 ( .A(learning_rate[9]), .Y(n23993) );
  AOI22XL U19666 ( .A0(n11536), .A1(data[9]), .B0(in_valid_d), .B1(w1[265]), 
        .Y(n9078) );
  INVXL U19667 ( .A(learning_rate[13]), .Y(n23990) );
  AOI22XL U19668 ( .A0(n4566), .A1(data[13]), .B0(in_valid_d), .B1(w1[269]), 
        .Y(n9079) );
  NAND2X1 U19669 ( .A(n9164), .B(target_temp[14]), .Y(n11529) );
  INVXL U19670 ( .A(n25157), .Y(n9081) );
  INVXL U19671 ( .A(learning_rate[5]), .Y(n23996) );
  AOI22XL U19672 ( .A0(n4566), .A1(data[5]), .B0(in_valid_d), .B1(w1[261]), 
        .Y(n9083) );
  AOI22X1 U19673 ( .A0(n4856), .A1(y12[10]), .B0(n14427), .B1(y10[10]), .Y(
        n9085) );
  INVXL U19674 ( .A(n25148), .Y(n9084) );
  INVXL U19675 ( .A(n25147), .Y(n9086) );
  AOI22XL U19676 ( .A0(n4566), .A1(data[12]), .B0(in_valid_d), .B1(w1[268]), 
        .Y(n9090) );
  INVXL U19677 ( .A(n25146), .Y(n9091) );
  INVXL U19678 ( .A(n24024), .Y(n9093) );
  INVX1 U19679 ( .A(learning_rate[0]), .Y(n24001) );
  AOI22XL U19680 ( .A0(n11536), .A1(data[0]), .B0(in_valid_d), .B1(w1[256]), 
        .Y(n9095) );
  NAND2X1 U19681 ( .A(n4826), .B(target_temp[0]), .Y(n11514) );
  AOI22XL U19682 ( .A0(n4566), .A1(data[2]), .B0(in_valid_d), .B1(w1[258]), 
        .Y(n9097) );
  NAND2X1 U19683 ( .A(n9164), .B(target_temp[2]), .Y(n11501) );
  OAI211X1 U19684 ( .A0(n24000), .A1(n25243), .B0(n9097), .C0(n11501), .Y(
        M2_b_2_) );
  AOI22XL U19685 ( .A0(n4856), .A1(y12[0]), .B0(n14427), .B1(y10[0]), .Y(n9099) );
  INVXL U19686 ( .A(n24266), .Y(n9098) );
  OAI211XL U19687 ( .A0(n25909), .A1(n9087), .B0(n9099), .C0(n9098), .Y(
        M2_a_0_) );
  AOI22XL U19688 ( .A0(n4566), .A1(data[17]), .B0(in_valid_d), .B1(w1[273]), 
        .Y(n9100) );
  INVXL U19689 ( .A(learning_rate[4]), .Y(n23998) );
  AOI22XL U19690 ( .A0(n4566), .A1(data[4]), .B0(in_valid_d), .B1(w1[260]), 
        .Y(n9102) );
  NAND2X1 U19691 ( .A(n4826), .B(target_temp[4]), .Y(n11508) );
  NOR2X1 U19692 ( .A(y10[31]), .B(n23973), .Y(n9108) );
  OAI22X4 U19693 ( .A0(n11057), .A1(n26218), .B0(n9107), .B1(n25950), .Y(
        n22867) );
  OAI22X1 U19694 ( .A0(n11057), .A1(n26219), .B0(n9107), .B1(n25892), .Y(
        n11159) );
  INVX1 U19695 ( .A(n11159), .Y(n26494) );
  OAI22X1 U19696 ( .A0(n11057), .A1(n26220), .B0(n9107), .B1(n25949), .Y(
        n11155) );
  OAI22X4 U19697 ( .A0(n11057), .A1(n26221), .B0(n9107), .B1(n25946), .Y(
        n23022) );
  CLKINVX3 U19698 ( .A(n26492), .Y(n26493) );
  CLKINVX3 U19699 ( .A(n11311), .Y(n23193) );
  OAI22X1 U19700 ( .A0(n23193), .A1(n26222), .B0(n9107), .B1(n25945), .Y(
        n11151) );
  INVX1 U19701 ( .A(n11151), .Y(n26491) );
  OAI22X1 U19702 ( .A0(n23193), .A1(n26223), .B0(n9107), .B1(n25944), .Y(
        n11147) );
  OAI22X1 U19703 ( .A0(n23193), .A1(n25993), .B0(n9107), .B1(n25890), .Y(
        n11141) );
  OAI22X4 U19704 ( .A0(n23193), .A1(n26230), .B0(n9107), .B1(n25939), .Y(
        n23089) );
  NOR2X1 U19705 ( .A(n9117), .B(n9116), .Y(n10676) );
  INVXL U19706 ( .A(learning_rate[29]), .Y(n21093) );
  INVXL U19707 ( .A(learning_rate[23]), .Y(n23065) );
  OAI21XL U19708 ( .A0(n9175), .A1(n9189), .B0(n9176), .Y(n9181) );
  OAI21XL U19709 ( .A0(n9174), .A1(n9170), .B0(n9171), .Y(n9168) );
  CMPR32X1 U19710 ( .A(n9169), .B(n10687), .C(n9168), .CO(n9184), .S(n24269)
         );
  CMPR32X1 U19711 ( .A(n9183), .B(n10686), .C(n9182), .CO(n9190), .S(n23661)
         );
  CMPR32X1 U19712 ( .A(n9185), .B(n10685), .C(n9184), .CO(n9182), .S(n24383)
         );
  CMPR32X1 U19713 ( .A(n9191), .B(n10684), .C(n9190), .CO(n20640), .S(n23662)
         );
  INVXL U19714 ( .A(n10287), .Y(n9196) );
  XNOR2X1 U19715 ( .A(M2_mult_x_15_n43), .B(n10342), .Y(n9230) );
  XNOR2X1 U19716 ( .A(M2_mult_x_15_n43), .B(n10341), .Y(n9209) );
  XOR2X1 U19717 ( .A(M2_a_2_), .B(M2_a_3_), .Y(n9199) );
  XNOR2X4 U19718 ( .A(M2_a_2_), .B(M2_mult_x_15_a_1_), .Y(n9906) );
  NAND2X2 U19719 ( .A(n9199), .B(n9906), .Y(n9445) );
  CLKBUFX8 U19720 ( .A(n9445), .Y(n9983) );
  INVX8 U19721 ( .A(n9907), .Y(n9904) );
  XOR2X1 U19722 ( .A(M2_a_4_), .B(M2_a_5_), .Y(n9200) );
  XNOR2X4 U19723 ( .A(M2_a_4_), .B(M2_a_3_), .Y(n9877) );
  NAND2X2 U19724 ( .A(n9200), .B(n9877), .Y(n9590) );
  XNOR2XL U19725 ( .A(M2_a_5_), .B(n10515), .Y(n9231) );
  XNOR2XL U19726 ( .A(M2_a_5_), .B(M2_mult_x_15_n1669), .Y(n9206) );
  OAI22XL U19727 ( .A0(n9979), .A1(n9231), .B0(n9877), .B1(n9206), .Y(n9245)
         );
  INVX8 U19728 ( .A(n9201), .Y(n9851) );
  XNOR2X1 U19729 ( .A(n10494), .B(n9836), .Y(n9240) );
  BUFX8 U19730 ( .A(M2_b_8_), .Y(n10312) );
  XNOR2X1 U19731 ( .A(n4808), .B(n10312), .Y(n9228) );
  OAI22XL U19732 ( .A0(n9504), .A1(n9228), .B0(n10496), .B1(n9208), .Y(n9242)
         );
  XNOR2X1 U19733 ( .A(n10339), .B(n10386), .Y(n9264) );
  BUFX8 U19734 ( .A(n10548), .Y(n10541) );
  XNOR2X1 U19735 ( .A(n25885), .B(n9836), .Y(n9210) );
  OAI22XL U19736 ( .A0(n10517), .A1(n9204), .B0(n10533), .B1(n9216), .Y(n9211)
         );
  XOR2X1 U19737 ( .A(M2_a_10_), .B(n21055), .Y(n9205) );
  OAI22XL U19738 ( .A0(n10325), .A1(n9226), .B0(n10326), .B1(n9272), .Y(n9282)
         );
  OAI22XL U19739 ( .A0(n9445), .A1(n9904), .B0(n9906), .B1(n9907), .Y(n9281)
         );
  XNOR2XL U19740 ( .A(n9886), .B(M2_mult_x_15_n1668), .Y(n9219) );
  OAI22XL U19741 ( .A0(n9979), .A1(n9206), .B0(n9877), .B1(n9219), .Y(n9280)
         );
  XNOR2XL U19742 ( .A(M2_a_7_), .B(n10515), .Y(n9220) );
  XNOR2X1 U19743 ( .A(M2_a_17_), .B(n10342), .Y(n9217) );
  XNOR2X1 U19744 ( .A(M2_mult_x_15_n43), .B(n10387), .Y(n9218) );
  XNOR2X1 U19745 ( .A(n25885), .B(n9839), .Y(n9360) );
  OAI22X1 U19746 ( .A0(n10541), .A1(n9210), .B0(n3174), .B1(n9360), .Y(n9364)
         );
  OAI2BB1XL U19747 ( .A0N(n9906), .A1N(n9983), .B0(n9904), .Y(n9363) );
  XNOR2X1 U19748 ( .A(n9841), .B(n10539), .Y(n9232) );
  XNOR2XL U19749 ( .A(n9841), .B(n10538), .Y(n9343) );
  OAI22XL U19750 ( .A0(n9966), .A1(n9232), .B0(n10159), .B1(n9343), .Y(n9355)
         );
  XNOR2XL U19751 ( .A(M2_a_17_), .B(n10341), .Y(n9340) );
  OAI22XL U19752 ( .A0(n9504), .A1(n9217), .B0(n10496), .B1(n9340), .Y(n9353)
         );
  XNOR2XL U19753 ( .A(n9851), .B(M2_mult_x_15_n1669), .Y(n9342) );
  OAI22XL U19754 ( .A0(n9551), .A1(n9220), .B0(n9838), .B1(n9342), .Y(n9337)
         );
  XNOR2XL U19755 ( .A(n9841), .B(n10335), .Y(n9223) );
  OAI21XL U19756 ( .A0(n3178), .A1(n9960), .B0(n10660), .Y(n9251) );
  XNOR2X1 U19757 ( .A(n9841), .B(n10514), .Y(n9233) );
  OAI22XL U19758 ( .A0(n9966), .A1(n9223), .B0(n10159), .B1(n9233), .Y(n9238)
         );
  OAI22X1 U19759 ( .A0(n10660), .A1(M2_b_2_), .B0(n3178), .B1(n9901), .Y(n9235) );
  BUFX8 U19760 ( .A(n10325), .Y(n10296) );
  XNOR2XL U19761 ( .A(n10324), .B(n10337), .Y(n9229) );
  OAI22XL U19762 ( .A0(n10296), .A1(n9229), .B0(n10326), .B1(n9226), .Y(n9234)
         );
  NAND2X2 U19763 ( .A(M2_mult_x_15_a_1_), .B(n9781), .Y(n9694) );
  XNOR2X1 U19764 ( .A(n25885), .B(n9892), .Y(n9302) );
  XNOR2X1 U19765 ( .A(n25885), .B(n9901), .Y(n9239) );
  XNOR2X1 U19766 ( .A(n10494), .B(n9874), .Y(n9318) );
  XNOR2X1 U19767 ( .A(n10494), .B(n9863), .Y(n9241) );
  OAI22XL U19768 ( .A0(n10517), .A1(n9318), .B0(n10533), .B1(n9241), .Y(n9303)
         );
  XNOR2X1 U19769 ( .A(n9851), .B(n10514), .Y(n9295) );
  XNOR2X1 U19770 ( .A(M2_a_17_), .B(n9839), .Y(n9296) );
  OAI22X1 U19771 ( .A0(n9504), .A1(n9296), .B0(n10496), .B1(n9228), .Y(n9262)
         );
  XNOR2X1 U19772 ( .A(n10324), .B(n10386), .Y(n9249) );
  OAI22XL U19773 ( .A0(n10296), .A1(n9249), .B0(n10326), .B1(n9229), .Y(n9261)
         );
  XNOR2XL U19774 ( .A(n9886), .B(n10538), .Y(n9254) );
  OAI22XL U19775 ( .A0(n9979), .A1(n9254), .B0(n9877), .B1(n9231), .Y(n9258)
         );
  OAI22XL U19776 ( .A0(n9966), .A1(n9233), .B0(n10159), .B1(n9232), .Y(n9275)
         );
  XNOR2X1 U19777 ( .A(n25885), .B(n9874), .Y(n9267) );
  OAI22X1 U19778 ( .A0(n10541), .A1(n9239), .B0(n3174), .B1(n9267), .Y(n9248)
         );
  OAI22XL U19779 ( .A0(n10517), .A1(n9241), .B0(n10533), .B1(n9240), .Y(n9247)
         );
  XNOR2XL U19780 ( .A(n9841), .B(n10337), .Y(n9322) );
  XNOR2X1 U19781 ( .A(n10324), .B(n10387), .Y(n9321) );
  OAI22X1 U19782 ( .A0(n10296), .A1(n9321), .B0(n10326), .B1(n9249), .Y(n9307)
         );
  XNOR2X1 U19783 ( .A(n10339), .B(n10342), .Y(n9381) );
  XNOR2X1 U19784 ( .A(M2_a_5_), .B(n10539), .Y(n9385) );
  OAI22XL U19785 ( .A0(n9979), .A1(n9385), .B0(n9877), .B1(n9254), .Y(n9376)
         );
  ADDFHX1 U19786 ( .A(n9257), .B(n9256), .CI(n9255), .CO(n9269), .S(n9374) );
  OAI22X1 U19787 ( .A0(n10541), .A1(n9267), .B0(n10329), .B1(n9266), .Y(n9276)
         );
  XNOR2X1 U19788 ( .A(n10324), .B(n10514), .Y(n9344) );
  OAI22XL U19789 ( .A0(n10296), .A1(n9272), .B0(n10326), .B1(n9344), .Y(n9358)
         );
  ADDFHX1 U19790 ( .A(n9277), .B(n9276), .CI(n9222), .CO(n9288), .S(n9283) );
  OAI22XL U19791 ( .A0(n9551), .A1(n9320), .B0(n9838), .B1(n9295), .Y(n9380)
         );
  XNOR2X1 U19792 ( .A(M2_a_17_), .B(n9836), .Y(n9319) );
  XNOR2X1 U19793 ( .A(M2_mult_x_15_n43), .B(n10312), .Y(n9317) );
  XNOR2XL U19794 ( .A(M2_mult_x_15_a_1_), .B(n23222), .Y(n9323) );
  OAI22X2 U19795 ( .A0(n9694), .A1(n9323), .B0(n9301), .B1(n3180), .Y(n9326)
         );
  XNOR2X1 U19796 ( .A(n10494), .B(n9901), .Y(n9398) );
  OAI22XL U19797 ( .A0(n9504), .A1(n9419), .B0(n10496), .B1(n9319), .Y(n9424)
         );
  BUFX3 U19798 ( .A(n10326), .Y(n9959) );
  XNOR2X1 U19799 ( .A(n9841), .B(n10386), .Y(n9420) );
  OAI22XL U19800 ( .A0(n9966), .A1(n9420), .B0(n10159), .B1(n9322), .Y(n9399)
         );
  XNOR2XL U19801 ( .A(M2_mult_x_15_a_1_), .B(n10515), .Y(n9405) );
  OAI22X1 U19802 ( .A0(n9963), .A1(n9405), .B0(n9323), .B1(n3180), .Y(n9404)
         );
  OAI22X1 U19803 ( .A0(n10541), .A1(n10540), .B0(n3174), .B1(n9324), .Y(n9403)
         );
  XNOR2X1 U19804 ( .A(n10339), .B(n10312), .Y(n9446) );
  XNOR2X1 U19805 ( .A(n9904), .B(n10539), .Y(n9444) );
  XNOR2XL U19806 ( .A(M2_a_5_), .B(n10335), .Y(n9439) );
  XNOR2X1 U19807 ( .A(M2_a_5_), .B(n10514), .Y(n9386) );
  OAI22XL U19808 ( .A0(n9979), .A1(n9439), .B0(n9877), .B1(n9386), .Y(n9447)
         );
  ADDFHX4 U19809 ( .A(n9330), .B(n9329), .CI(n9328), .CO(n9268), .S(n9370) );
  XNOR2X1 U19810 ( .A(M2_a_17_), .B(n10387), .Y(n9460) );
  XNOR2XL U19811 ( .A(n9851), .B(n9341), .Y(n9479) );
  OAI22XL U19812 ( .A0(n9551), .A1(n9342), .B0(n9838), .B1(n9479), .Y(n9469)
         );
  XNOR2XL U19813 ( .A(n9841), .B(n10515), .Y(n9463) );
  OAI22XL U19814 ( .A0(n9966), .A1(n9343), .B0(n10159), .B1(n9463), .Y(n9468)
         );
  XNOR2X1 U19815 ( .A(n10324), .B(n10539), .Y(n9459) );
  OAI22XL U19816 ( .A0(n10296), .A1(n9344), .B0(n10326), .B1(n9459), .Y(n9482)
         );
  XNOR2XL U19817 ( .A(n10339), .B(n10335), .Y(n9461) );
  OAI22XL U19818 ( .A0(n10368), .A1(n9345), .B0(n10369), .B1(n9461), .Y(n9481)
         );
  CMPR32X1 U19819 ( .A(n3182), .B(n9901), .C(n9346), .CO(n9480), .S(n9356) );
  CMPR32X1 U19820 ( .A(n9355), .B(n9354), .C(n9353), .CO(n9458), .S(n9332) );
  INVXL U19821 ( .A(n9874), .Y(n9467) );
  OAI22XL U19822 ( .A0(n9979), .A1(n9886), .B0(n9877), .B1(n9878), .Y(n9465)
         );
  XNOR2X1 U19823 ( .A(n25885), .B(n10312), .Y(n9462) );
  OAI22XL U19824 ( .A0(n10517), .A1(n9362), .B0(n10533), .B1(n9464), .Y(n9477)
         );
  OAI22XL U19825 ( .A0(n9979), .A1(n9386), .B0(n9877), .B1(n9385), .Y(n9422)
         );
  ADDFHX1 U19826 ( .A(n9392), .B(n9391), .CI(n9390), .CO(n9387), .S(n10064) );
  XNOR2X1 U19827 ( .A(n25885), .B(n9960), .Y(n9397) );
  OAI22XL U19828 ( .A0(n10548), .A1(n9397), .B0(n3174), .B1(n9396), .Y(n9451)
         );
  XNOR2X1 U19829 ( .A(n10494), .B(n9892), .Y(n9406) );
  OAI22XL U19830 ( .A0(n10517), .A1(n9406), .B0(n10533), .B1(n9398), .Y(n9450)
         );
  XNOR2X1 U19831 ( .A(M2_mult_x_15_n43), .B(n9836), .Y(n9435) );
  CMPR22X1 U19832 ( .A(n9404), .B(n9403), .CO(n9432), .S(n10075) );
  NOR2BX1 U19833 ( .AN(n9960), .B(n3174), .Y(n9598) );
  XNOR2XL U19834 ( .A(M2_mult_x_15_a_1_), .B(n10538), .Y(n9441) );
  XNOR2X1 U19835 ( .A(M2_a_17_), .B(n9874), .Y(n9434) );
  XNOR2X1 U19836 ( .A(n9841), .B(n10387), .Y(n9443) );
  XNOR2XL U19837 ( .A(n9851), .B(n10337), .Y(n9440) );
  OAI22XL U19838 ( .A0(n9551), .A1(n9440), .B0(n9838), .B1(n9421), .Y(n9436)
         );
  CMPR32X1 U19839 ( .A(n9426), .B(n9425), .C(n9424), .CO(n9429), .S(n10068) );
  XNOR2X1 U19840 ( .A(M2_a_17_), .B(n9901), .Y(n9602) );
  OAI22X1 U19841 ( .A0(n9504), .A1(n9602), .B0(n10496), .B1(n9434), .Y(n9622)
         );
  XNOR2X1 U19842 ( .A(M2_mult_x_15_n43), .B(n9863), .Y(n9616) );
  ADDFHX1 U19843 ( .A(n9438), .B(n9437), .CI(n9436), .CO(n10070), .S(n10091)
         );
  XNOR2XL U19844 ( .A(M2_a_5_), .B(M2_b_15_), .Y(n9589) );
  XNOR2X1 U19845 ( .A(n9851), .B(n10386), .Y(n9592) );
  OAI22XL U19846 ( .A0(n9551), .A1(n9592), .B0(n9838), .B1(n9440), .Y(n9625)
         );
  XNOR2X1 U19847 ( .A(M2_mult_x_15_a_1_), .B(n10539), .Y(n9595) );
  XNOR2X1 U19848 ( .A(n9904), .B(n10514), .Y(n9614) );
  XNOR2X1 U19849 ( .A(n10339), .B(n9839), .Y(n9591) );
  OAI22XL U19850 ( .A0(n10368), .A1(n9591), .B0(n9780), .B1(n9446), .Y(n9604)
         );
  CMPR32X1 U19851 ( .A(n9452), .B(n9451), .C(n9450), .CO(n10073), .S(n10087)
         );
  CMPR32X1 U19852 ( .A(n9455), .B(n9454), .C(n9453), .CO(n9491), .S(n9488) );
  XNOR2XL U19853 ( .A(n10324), .B(n10538), .Y(n9516) );
  XNOR2X1 U19854 ( .A(n10339), .B(n10514), .Y(n9503) );
  OAI22XL U19855 ( .A0(n10368), .A1(n9461), .B0(n10369), .B1(n9503), .Y(n9513)
         );
  XNOR2XL U19856 ( .A(n9841), .B(M2_mult_x_15_n1669), .Y(n9501) );
  OAI22XL U19857 ( .A0(n10517), .A1(n9464), .B0(n10533), .B1(n9507), .Y(n9510)
         );
  OAI22XL U19858 ( .A0(n10660), .A1(n9836), .B0(n10659), .B1(n9839), .Y(n9517)
         );
  CMPR32X1 U19859 ( .A(n9470), .B(n9469), .C(n9468), .CO(n9492), .S(n9475) );
  OAI22XL U19860 ( .A0(n9551), .A1(n9479), .B0(n9838), .B1(n9851), .Y(n9499)
         );
  OAI2BB1XL U19861 ( .A0N(n9877), .A1N(n9590), .B0(M2_a_5_), .Y(n9498) );
  CMPR32X1 U19862 ( .A(n9482), .B(n9481), .C(n9480), .CO(n9495), .S(n9474) );
  XNOR2XL U19863 ( .A(n9841), .B(M2_mult_x_15_n1668), .Y(n9550) );
  OAI22XL U19864 ( .A0(n4570), .A1(n9502), .B0(n10403), .B1(n9549), .Y(n9534)
         );
  XNOR2X1 U19865 ( .A(n10339), .B(n10539), .Y(n9543) );
  OAI22XL U19866 ( .A0(n10368), .A1(n9503), .B0(n10369), .B1(n9543), .Y(n9533)
         );
  XNOR2XL U19867 ( .A(M2_a_17_), .B(n10337), .Y(n9538) );
  OAI22XL U19868 ( .A0(n9504), .A1(n9505), .B0(n10496), .B1(n9538), .Y(n9548)
         );
  XNOR2X1 U19869 ( .A(n25885), .B(n10342), .Y(n9536) );
  OAI22X1 U19870 ( .A0(n10541), .A1(n9506), .B0(n10329), .B1(n9536), .Y(n9547)
         );
  XNOR2X1 U19871 ( .A(n10494), .B(n10387), .Y(n9537) );
  OAI22XL U19872 ( .A0(n10517), .A1(n9507), .B0(n10533), .B1(n9537), .Y(n9546)
         );
  CMPR32X1 U19873 ( .A(n9512), .B(n9511), .C(n9510), .CO(n9532), .S(n9519) );
  XNOR2XL U19874 ( .A(n10324), .B(n10515), .Y(n9542) );
  OAI22XL U19875 ( .A0(n10296), .A1(n9516), .B0(n10326), .B1(n9542), .Y(n9541)
         );
  CMPR32X1 U19876 ( .A(n9874), .B(n9863), .C(n9517), .CO(n9540), .S(n9494) );
  OAI22XL U19877 ( .A0(n9551), .A1(n9851), .B0(n9838), .B1(n9201), .Y(n9544)
         );
  CMPR32X1 U19878 ( .A(n9526), .B(n9525), .C(n9524), .CO(n9560), .S(n9557) );
  XNOR2XL U19879 ( .A(n25885), .B(n10341), .Y(n9580) );
  XNOR2XL U19880 ( .A(M2_a_17_), .B(M2_b_15_), .Y(n9573) );
  OAI22XL U19881 ( .A0(n9504), .A1(n9538), .B0(n10496), .B1(n9573), .Y(n9570)
         );
  XNOR2XL U19882 ( .A(n10324), .B(M2_mult_x_15_n1669), .Y(n9574) );
  OAI22XL U19883 ( .A0(n10296), .A1(n9542), .B0(n10326), .B1(n9574), .Y(n9578)
         );
  XNOR2X1 U19884 ( .A(n10339), .B(n10538), .Y(n9575) );
  OAI22XL U19885 ( .A0(n10368), .A1(n9543), .B0(n10369), .B1(n9575), .Y(n9577)
         );
  OAI22XL U19886 ( .A0(n10660), .A1(n10312), .B0(n3178), .B1(n10311), .Y(n9582) );
  XNOR2X1 U19887 ( .A(M2_mult_x_15_n43), .B(n10514), .Y(n9579) );
  OAI2BB1XL U19888 ( .A0N(n9838), .A1N(n9551), .B0(M2_a_7_), .Y(n9583) );
  ADDFHX1 U19889 ( .A(n9563), .B(n9562), .CI(n9561), .CO(n10147), .S(n9564) );
  ADDFHX1 U19890 ( .A(n9572), .B(n9571), .CI(n9570), .CO(n10153), .S(n9568) );
  XNOR2XL U19891 ( .A(M2_a_17_), .B(n10335), .Y(n10157) );
  XNOR2XL U19892 ( .A(n10339), .B(n10515), .Y(n10160) );
  OAI22XL U19893 ( .A0(n10368), .A1(n9575), .B0(n10369), .B1(n10160), .Y(
        n10154) );
  CMPR32X1 U19894 ( .A(n9578), .B(n9577), .C(n9576), .CO(n10151), .S(n9563) );
  XNOR2X1 U19895 ( .A(M2_mult_x_15_n43), .B(n10539), .Y(n10169) );
  XNOR2X1 U19896 ( .A(n25885), .B(n10387), .Y(n10161) );
  XNOR2XL U19897 ( .A(n10494), .B(n10337), .Y(n10162) );
  CMPR32X1 U19898 ( .A(n9836), .B(n9839), .C(n9582), .CO(n10168), .S(n9576) );
  OAI22XL U19899 ( .A0(n9966), .A1(n9841), .B0(n10159), .B1(n9843), .Y(n10170)
         );
  ADDFHX1 U19900 ( .A(n9585), .B(n9584), .CI(n9583), .CO(n10166), .S(n9586) );
  ADDFHX1 U19901 ( .A(n9588), .B(n9587), .CI(n9586), .CO(n10148), .S(n9562) );
  XNOR2XL U19902 ( .A(M2_a_5_), .B(n10337), .Y(n9607) );
  OAI22XL U19903 ( .A0(n9590), .A1(n9607), .B0(n9877), .B1(n9589), .Y(n9629)
         );
  XNOR2X1 U19904 ( .A(n10339), .B(n9836), .Y(n9608) );
  OAI22XL U19905 ( .A0(n10368), .A1(n9608), .B0(n9780), .B1(n9591), .Y(n9628)
         );
  OAI22XL U19906 ( .A0(n9551), .A1(n9630), .B0(n9838), .B1(n9592), .Y(n9627)
         );
  CMPR22X1 U19907 ( .A(n9594), .B(n9593), .CO(n9624), .S(n9638) );
  NOR2BX1 U19908 ( .AN(n9960), .B(n10533), .Y(n9635) );
  XNOR2X1 U19909 ( .A(M2_a_17_), .B(n9892), .Y(n9603) );
  XNOR2X1 U19910 ( .A(n10324), .B(n9839), .Y(n9639) );
  XNOR2X1 U19911 ( .A(n10324), .B(n10312), .Y(n9601) );
  OAI22XL U19912 ( .A0(n10296), .A1(n9639), .B0(n9959), .B1(n9601), .Y(n9647)
         );
  XNOR2X1 U19913 ( .A(M2_mult_x_15_n43), .B(n9874), .Y(n9617) );
  XNOR2XL U19914 ( .A(n9904), .B(n10335), .Y(n9615) );
  OAI22XL U19915 ( .A0(n9983), .A1(n9640), .B0(n9906), .B1(n9615), .Y(n9645)
         );
  ADDFHX1 U19916 ( .A(n9598), .B(n9597), .CI(n9596), .CO(n10074), .S(n10079)
         );
  OAI22X1 U19917 ( .A0(n10296), .A1(n9601), .B0(n9959), .B1(n9600), .Y(n9610)
         );
  OAI22XL U19918 ( .A0(n9504), .A1(n9603), .B0(n10496), .B1(n9602), .Y(n9609)
         );
  XNOR2X1 U19919 ( .A(n9841), .B(n10311), .Y(n9656) );
  XNOR2X1 U19920 ( .A(n9841), .B(M2_b_10_), .Y(n9613) );
  OAI22XL U19921 ( .A0(n9966), .A1(n9656), .B0(n10159), .B1(n9613), .Y(n9644)
         );
  XNOR2X1 U19922 ( .A(n9886), .B(n10386), .Y(n9641) );
  BUFX3 U19923 ( .A(n9877), .Y(n9977) );
  OAI22X1 U19924 ( .A0(n9590), .A1(n9641), .B0(n9877), .B1(n9607), .Y(n9643)
         );
  XNOR2X1 U19925 ( .A(n10339), .B(n9863), .Y(n9654) );
  OAI22XL U19926 ( .A0(n10368), .A1(n9654), .B0(n9780), .B1(n9608), .Y(n9642)
         );
  OAI22XL U19927 ( .A0(n9966), .A1(n9613), .B0(n10159), .B1(n9612), .Y(n9620)
         );
  OAI22X1 U19928 ( .A0(n9983), .A1(n9615), .B0(n9906), .B1(n9614), .Y(n9619)
         );
  ADDFHX1 U19929 ( .A(n9623), .B(n9622), .CI(n9621), .CO(n10092), .S(n10081)
         );
  CMPR32X1 U19930 ( .A(n9626), .B(n9625), .C(n9624), .CO(n10090), .S(n10080)
         );
  CMPR32X1 U19931 ( .A(n9629), .B(n9628), .C(n9627), .CO(n10095), .S(n9664) );
  OAI22XL U19932 ( .A0(n9551), .A1(n9655), .B0(n9974), .B1(n9630), .Y(n9661)
         );
  XNOR2X1 U19933 ( .A(M2_mult_x_15_a_1_), .B(n10335), .Y(n9665) );
  ADDFHX1 U19934 ( .A(n9635), .B(n9634), .CI(n9633), .CO(n9637), .S(n9659) );
  XNOR2X1 U19935 ( .A(n10324), .B(n9836), .Y(n9674) );
  OAI22XL U19936 ( .A0(n10325), .A1(n9674), .B0(n9959), .B1(n9639), .Y(n9672)
         );
  XNOR2XL U19937 ( .A(M2_a_3_), .B(n10337), .Y(n9668) );
  BUFX3 U19938 ( .A(n9906), .Y(n9981) );
  XNOR2X1 U19939 ( .A(n9886), .B(n10387), .Y(n9673) );
  OAI22XL U19940 ( .A0(n9979), .A1(n9673), .B0(n9877), .B1(n9641), .Y(n9670)
         );
  ADDFHX1 U19941 ( .A(n9647), .B(n9646), .CI(n9645), .CO(n9636), .S(n9681) );
  XNOR2X1 U19942 ( .A(M2_mult_x_15_n43), .B(n9892), .Y(n9666) );
  XNOR2X1 U19943 ( .A(n10339), .B(n9874), .Y(n9669) );
  XNOR2X1 U19944 ( .A(n9851), .B(n10342), .Y(n9675) );
  OAI22XL U19945 ( .A0(n9551), .A1(n9675), .B0(n9974), .B1(n9655), .Y(n9680)
         );
  XNOR2X1 U19946 ( .A(n9841), .B(n10312), .Y(n9667) );
  OAI22XL U19947 ( .A0(n9966), .A1(n9667), .B0(n10159), .B1(n9656), .Y(n9679)
         );
  ADDFHX1 U19948 ( .A(n9664), .B(n9663), .CI(n9662), .CO(n10105), .S(n9689) );
  OAI22X2 U19949 ( .A0(n9694), .A1(n9693), .B0(n9665), .B1(n3180), .Y(n9697)
         );
  XNOR2XL U19950 ( .A(M2_mult_x_15_n43), .B(n3182), .Y(n9700) );
  XNOR2X1 U19951 ( .A(n9841), .B(n9839), .Y(n9699) );
  XNOR2X1 U19952 ( .A(n10339), .B(n9901), .Y(n9702) );
  OAI22XL U19953 ( .A0(n10368), .A1(n9702), .B0(n9780), .B1(n9669), .Y(n9709)
         );
  ADDFHX1 U19954 ( .A(n9672), .B(n9671), .CI(n9670), .CO(n9683), .S(n9703) );
  XNOR2XL U19955 ( .A(n9886), .B(n10341), .Y(n9721) );
  OAI22X1 U19956 ( .A0(n10296), .A1(n9707), .B0(n9959), .B1(n9674), .Y(n9713)
         );
  OAI22XL U19957 ( .A0(n9551), .A1(n9708), .B0(n9974), .B1(n9675), .Y(n9712)
         );
  CMPR32X1 U19958 ( .A(n9680), .B(n9679), .C(n9678), .CO(n9691), .S(n9718) );
  ADDFHX1 U19959 ( .A(n9683), .B(n9682), .CI(n9681), .CO(n9686), .S(n9715) );
  XNOR2XL U19960 ( .A(M2_mult_x_15_a_1_), .B(n10337), .Y(n9723) );
  XNOR2X1 U19961 ( .A(n9841), .B(n9836), .Y(n9728) );
  XNOR2X1 U19962 ( .A(M2_mult_x_15_n43), .B(n9960), .Y(n9701) );
  XNOR2X1 U19963 ( .A(n10339), .B(n9892), .Y(n9724) );
  OAI22XL U19964 ( .A0(n10368), .A1(n9724), .B0(n9780), .B1(n9702), .Y(n9731)
         );
  XNOR2X1 U19965 ( .A(n9904), .B(n10387), .Y(n9730) );
  XNOR2X1 U19966 ( .A(n10324), .B(n9874), .Y(n9729) );
  OAI22X1 U19967 ( .A0(n10296), .A1(n9729), .B0(n9959), .B1(n9707), .Y(n9745)
         );
  XNOR2X1 U19968 ( .A(n9851), .B(n10312), .Y(n9735) );
  OAI22XL U19969 ( .A0(n9551), .A1(n9735), .B0(n9974), .B1(n9708), .Y(n9744)
         );
  ADDFHX1 U19970 ( .A(n9711), .B(n9710), .CI(n9709), .CO(n9704), .S(n9742) );
  XNOR2X1 U19971 ( .A(n9886), .B(n10342), .Y(n9734) );
  OAI22XL U19972 ( .A0(n9979), .A1(n9734), .B0(n9977), .B1(n9721), .Y(n9749)
         );
  OAI22X1 U19973 ( .A0(n9963), .A1(n9736), .B0(n9723), .B1(n3180), .Y(n9751)
         );
  XNOR2X1 U19974 ( .A(n10339), .B(n3182), .Y(n9772) );
  OAI22XL U19975 ( .A0(n10368), .A1(n9772), .B0(n9780), .B1(n9724), .Y(n9750)
         );
  OAI22XL U19976 ( .A0(n9983), .A1(n9754), .B0(n9981), .B1(n9730), .Y(n9756)
         );
  XNOR2X1 U19977 ( .A(n9886), .B(n10311), .Y(n9755) );
  XNOR2X1 U19978 ( .A(M2_mult_x_15_a_1_), .B(n10387), .Y(n9782) );
  OAI22XL U19979 ( .A0(n10368), .A1(n10338), .B0(n10369), .B1(n9737), .Y(n9778) );
  ADDFHX1 U19980 ( .A(n9746), .B(n9745), .CI(n9744), .CO(n9743), .S(n9789) );
  XNOR2X1 U19981 ( .A(n9841), .B(n9874), .Y(n9798) );
  XNOR2X1 U19982 ( .A(n9886), .B(n10312), .Y(n9786) );
  CMPR32X1 U19983 ( .A(n9761), .B(n9760), .C(n9759), .CO(n9766), .S(n9827) );
  XNOR2X1 U19984 ( .A(n9851), .B(n9836), .Y(n9784) );
  OAI22XL U19985 ( .A0(n9551), .A1(n9784), .B0(n9974), .B1(n9771), .Y(n9795)
         );
  XNOR2X1 U19986 ( .A(n10339), .B(n9960), .Y(n9773) );
  XNOR2X1 U19987 ( .A(n10324), .B(n9892), .Y(n9783) );
  OAI22XL U19988 ( .A0(n10296), .A1(n9783), .B0(n9959), .B1(n9774), .Y(n9793)
         );
  ADDHXL U19989 ( .A(n9779), .B(n9778), .CO(n9775), .S(n9811) );
  XNOR2XL U19990 ( .A(n10324), .B(n3182), .Y(n9813) );
  OAI22XL U19991 ( .A0(n10296), .A1(n9813), .B0(n9959), .B1(n9783), .Y(n9800)
         );
  XNOR2X1 U19992 ( .A(n9851), .B(n9863), .Y(n9812) );
  OAI22XL U19993 ( .A0(n9551), .A1(n9812), .B0(n9974), .B1(n9784), .Y(n9822)
         );
  XNOR2X1 U19994 ( .A(n9886), .B(n9839), .Y(n9816) );
  OAI22XL U19995 ( .A0(n9979), .A1(n9816), .B0(n9977), .B1(n9786), .Y(n9820)
         );
  CMPR32X1 U19996 ( .A(n9795), .B(n9794), .C(n9793), .CO(n9805), .S(n9825) );
  XNOR2X1 U19997 ( .A(n9841), .B(n9901), .Y(n9817) );
  XNOR2X1 U19998 ( .A(M2_mult_x_15_a_1_), .B(M2_b_10_), .Y(n9961) );
  ADDFHX1 U19999 ( .A(n9811), .B(n9810), .CI(n9809), .CO(n9803), .S(n10016) );
  XNOR2X1 U20000 ( .A(n9851), .B(n9874), .Y(n9973) );
  OAI22XL U20001 ( .A0(n9551), .A1(n9973), .B0(n9974), .B1(n9812), .Y(n9986)
         );
  XNOR2X1 U20002 ( .A(n10324), .B(n9960), .Y(n9814) );
  OAI22XL U20003 ( .A0(n10296), .A1(n9814), .B0(n9959), .B1(n9813), .Y(n9985)
         );
  OAI22XL U20004 ( .A0(n9983), .A1(n9980), .B0(n9981), .B1(n9815), .Y(n9984)
         );
  OAI22XL U20005 ( .A0(n9979), .A1(n9976), .B0(n9977), .B1(n9816), .Y(n9956)
         );
  XNOR2X1 U20006 ( .A(n9841), .B(n9892), .Y(n9964) );
  CMPR22X1 U20007 ( .A(n9819), .B(n9818), .CO(n10018), .S(n9954) );
  NOR2XL U20008 ( .A(n10043), .B(n10042), .Y(n9826) );
  NOR2XL U20009 ( .A(n10046), .B(n9826), .Y(n9833) );
  NOR2X1 U20010 ( .A(n10048), .B(n10047), .Y(n9832) );
  XNOR2X1 U20011 ( .A(n9851), .B(n9892), .Y(n9846) );
  XNOR2X1 U20012 ( .A(n9851), .B(n9901), .Y(n9975) );
  OAI22XL U20013 ( .A0(n9551), .A1(n9846), .B0(n9974), .B1(n9975), .Y(n9969)
         );
  XNOR2XL U20014 ( .A(n9841), .B(n3182), .Y(n9965) );
  XNOR2X1 U20015 ( .A(n9886), .B(n9874), .Y(n9835) );
  XNOR2X1 U20016 ( .A(n9886), .B(n9863), .Y(n9978) );
  OAI22XL U20017 ( .A0(n9979), .A1(n9835), .B0(n9977), .B1(n9978), .Y(n9967)
         );
  XNOR2X1 U20018 ( .A(n9904), .B(n9863), .Y(n9850) );
  OAI22XL U20019 ( .A0(n9983), .A1(n9850), .B0(n9981), .B1(n9840), .Y(n9857)
         );
  XNOR2X1 U20020 ( .A(n9886), .B(n9901), .Y(n9854) );
  OAI22XL U20021 ( .A0(n9979), .A1(n9854), .B0(n9977), .B1(n9835), .Y(n9856)
         );
  XNOR2X1 U20022 ( .A(M2_mult_x_15_a_1_), .B(n9836), .Y(n9864) );
  XNOR2X1 U20023 ( .A(M2_mult_x_15_a_1_), .B(n9839), .Y(n9845) );
  OAI22XL U20024 ( .A0(n9963), .A1(n9864), .B0(n9845), .B1(n3180), .Y(n9862)
         );
  NAND2BXL U20025 ( .AN(n9960), .B(n9851), .Y(n9837) );
  OAI22XL U20026 ( .A0(n9551), .A1(n9201), .B0(n9838), .B1(n9837), .Y(n9861)
         );
  OAI22XL U20027 ( .A0(n9983), .A1(n9840), .B0(n9981), .B1(n9982), .Y(n9992)
         );
  NAND2BXL U20028 ( .AN(n9960), .B(n9841), .Y(n9842) );
  OAI22XL U20029 ( .A0(n9966), .A1(n9843), .B0(n10159), .B1(n9842), .Y(n9957)
         );
  XNOR2XL U20030 ( .A(n9851), .B(n3182), .Y(n9852) );
  OAI22XL U20031 ( .A0(n9551), .A1(n9852), .B0(n9974), .B1(n9846), .Y(n9847)
         );
  OAI22XL U20032 ( .A0(n9983), .A1(n9873), .B0(n9981), .B1(n9850), .Y(n9868)
         );
  OAI22XL U20033 ( .A0(n9551), .A1(n9853), .B0(n9974), .B1(n9852), .Y(n9867)
         );
  XNOR2X1 U20034 ( .A(n9886), .B(n9892), .Y(n9865) );
  NOR2XL U20035 ( .A(n9947), .B(n9946), .Y(n9950) );
  CMPR32X1 U20036 ( .A(n9860), .B(n9859), .C(n9858), .CO(n9946), .S(n9945) );
  ADDHXL U20037 ( .A(n9862), .B(n9861), .CO(n9855), .S(n9872) );
  NOR2BX1 U20038 ( .AN(n9960), .B(n9974), .Y(n9881) );
  XNOR2X1 U20039 ( .A(M2_mult_x_15_a_1_), .B(n9863), .Y(n9875) );
  XNOR2X1 U20040 ( .A(n9886), .B(n3182), .Y(n9887) );
  CMPR32X1 U20041 ( .A(n9868), .B(n9867), .C(n9866), .CO(n9859), .S(n9870) );
  NOR2XL U20042 ( .A(n9945), .B(n9944), .Y(n9869) );
  NOR2XL U20043 ( .A(n9950), .B(n9869), .Y(n9953) );
  XNOR2X1 U20044 ( .A(M2_mult_x_15_a_1_), .B(n9874), .Y(n9912) );
  OAI22XL U20045 ( .A0(n9963), .A1(n9912), .B0(n9875), .B1(n3180), .Y(n9890)
         );
  OR2X2 U20046 ( .A(n9937), .B(n9936), .Y(n9940) );
  ADDHXL U20047 ( .A(n9890), .B(n9889), .CO(n9883), .S(n9923) );
  OR2X2 U20048 ( .A(n9935), .B(n9934), .Y(n9891) );
  NAND2XL U20049 ( .A(n9940), .B(n9891), .Y(n9943) );
  INVXL U20050 ( .A(n9897), .Y(n9900) );
  INVXL U20051 ( .A(n9893), .Y(n9894) );
  NAND2XL U20052 ( .A(n9895), .B(n9894), .Y(n9899) );
  NAND2XL U20053 ( .A(n9897), .B(n9896), .Y(n9898) );
  OAI21XL U20054 ( .A0(n9900), .A1(n9899), .B0(n9898), .Y(n9911) );
  XNOR2X1 U20055 ( .A(M2_mult_x_15_a_1_), .B(n9901), .Y(n9913) );
  XNOR2X1 U20056 ( .A(n9904), .B(n3182), .Y(n9915) );
  AOI21XL U20057 ( .A0(n9911), .A1(n9908), .B0(n6201), .Y(n9922) );
  NOR2BXL U20058 ( .AN(n9960), .B(n9977), .Y(n9928) );
  NOR2XL U20059 ( .A(n9919), .B(n9918), .Y(n9921) );
  NAND2XL U20060 ( .A(n9919), .B(n9918), .Y(n9920) );
  OAI21XL U20061 ( .A0(n9922), .A1(n9921), .B0(n9920), .Y(n9933) );
  CMPR32X1 U20062 ( .A(n9925), .B(n9924), .C(n9923), .CO(n9934), .S(n9931) );
  CMPR32X1 U20063 ( .A(n9928), .B(n9927), .C(n9926), .CO(n9930), .S(n9919) );
  AND2X2 U20064 ( .A(n9935), .B(n9934), .Y(n9939) );
  AOI21XL U20065 ( .A0(n9940), .A1(n9939), .B0(n9938), .Y(n9941) );
  OAI21XL U20066 ( .A0(n9943), .A1(n9942), .B0(n9941), .Y(n9952) );
  NAND2XL U20067 ( .A(n9945), .B(n9944), .Y(n9949) );
  NAND2XL U20068 ( .A(n9947), .B(n9946), .Y(n9948) );
  OAI21XL U20069 ( .A0(n9950), .A1(n9949), .B0(n9948), .Y(n9951) );
  AOI21XL U20070 ( .A0(n9953), .A1(n9952), .B0(n9951), .Y(n10013) );
  CMPR32X1 U20071 ( .A(n9956), .B(n9955), .C(n9954), .CO(n10024), .S(n10031)
         );
  NOR2BX1 U20072 ( .AN(n9960), .B(n9959), .Y(n9972) );
  OAI22XL U20073 ( .A0(n9966), .A1(n9965), .B0(n10159), .B1(n9964), .Y(n9970)
         );
  CMPR32X1 U20074 ( .A(n9972), .B(n9971), .C(n9970), .CO(n10022), .S(n9994) );
  OAI22XL U20075 ( .A0(n9551), .A1(n9975), .B0(n9974), .B1(n9973), .Y(n9989)
         );
  OAI22XL U20076 ( .A0(n9983), .A1(n9982), .B0(n9981), .B1(n9980), .Y(n9987)
         );
  CMPR32X1 U20077 ( .A(n9986), .B(n9985), .C(n9984), .CO(n10025), .S(n10020)
         );
  CMPR32X1 U20078 ( .A(n9989), .B(n9988), .C(n9987), .CO(n10021), .S(n9999) );
  ADDFHX1 U20079 ( .A(n9992), .B(n9991), .CI(n9990), .CO(n9998), .S(n10000) );
  NOR2XL U20080 ( .A(n10007), .B(n10006), .Y(n9996) );
  INVXL U20081 ( .A(n9996), .Y(n10010) );
  CMPR32X1 U20082 ( .A(n9999), .B(n9998), .C(n9997), .CO(n10006), .S(n10005)
         );
  CMPR32X1 U20083 ( .A(n10002), .B(n10001), .C(n10000), .CO(n10004), .S(n9947)
         );
  NAND2XL U20084 ( .A(n10003), .B(n10010), .Y(n10012) );
  AND2X2 U20085 ( .A(n10007), .B(n10006), .Y(n10008) );
  AOI21XL U20086 ( .A0(n10010), .A1(n10009), .B0(n10008), .Y(n10011) );
  OAI21XL U20087 ( .A0(n10013), .A1(n10012), .B0(n10011), .Y(n10041) );
  CMPR32X1 U20088 ( .A(n10019), .B(n10018), .C(n10017), .CO(n9823), .S(n10028)
         );
  CMPR32X1 U20089 ( .A(n10028), .B(n10027), .C(n10026), .CO(n10035), .S(n10034) );
  NOR2XL U20090 ( .A(n10034), .B(n10033), .Y(n10032) );
  NAND2XL U20091 ( .A(n10034), .B(n10033), .Y(n10038) );
  NAND2XL U20092 ( .A(n10036), .B(n10035), .Y(n10037) );
  AND2X2 U20093 ( .A(n10048), .B(n10047), .Y(n10049) );
  ADDFHX4 U20094 ( .A(n10061), .B(n10060), .CI(n10059), .CO(n10128), .S(n10124) );
  CMPR32X1 U20095 ( .A(n10076), .B(n10075), .C(n10074), .CO(n10071), .S(n10104) );
  ADDFHX1 U20096 ( .A(n10089), .B(n10088), .CI(n10087), .CO(n10084), .S(n10110) );
  ADDFHX1 U20097 ( .A(n10095), .B(n10094), .CI(n10093), .CO(n10108), .S(n10116) );
  OAI22XL U20098 ( .A0(n10325), .A1(n10158), .B0(n10326), .B1(n10324), .Y(
        n10298) );
  XNOR2XL U20099 ( .A(n10339), .B(M2_mult_x_15_n1669), .Y(n10308) );
  OAI22XL U20100 ( .A0(n10368), .A1(n10160), .B0(n10369), .B1(n10308), .Y(
        n10307) );
  XNOR2XL U20101 ( .A(n10494), .B(M2_b_15_), .Y(n10299) );
  OAI22XL U20102 ( .A0(n10532), .A1(n10162), .B0(n10533), .B1(n10299), .Y(
        n10305) );
  XNOR2X1 U20103 ( .A(M2_mult_x_15_n43), .B(n10538), .Y(n10309) );
  OAI22XL U20104 ( .A0(n10660), .A1(n10342), .B0(n3178), .B1(n10341), .Y(
        n10310) );
  CMPR32X1 U20105 ( .A(n10174), .B(n10173), .C(n10172), .CO(n10289), .S(n10145) );
  INVXL U20106 ( .A(n10446), .Y(n10177) );
  NAND2X2 U20107 ( .A(n10176), .B(n10175), .Y(n10464) );
  INVXL U20108 ( .A(n10179), .Y(n10229) );
  INVXL U20109 ( .A(n10180), .Y(n10224) );
  NAND2XL U20110 ( .A(n10229), .B(n10224), .Y(n10185) );
  INVXL U20111 ( .A(n10223), .Y(n10183) );
  INVXL U20112 ( .A(n10186), .Y(n10188) );
  INVXL U20113 ( .A(n10228), .Y(n10192) );
  NAND2XL U20114 ( .A(n10229), .B(n10192), .Y(n10194) );
  INVXL U20115 ( .A(n10191), .Y(n10231) );
  INVXL U20116 ( .A(n10201), .Y(n10203) );
  INVXL U20117 ( .A(n10218), .Y(n10204) );
  NAND2X1 U20118 ( .A(n10204), .B(n10217), .Y(n10205) );
  XOR2X2 U20119 ( .A(n10243), .B(n10205), .Y(n19073) );
  NAND2XL U20120 ( .A(n10240), .B(n10245), .Y(n10212) );
  INVXL U20121 ( .A(n10244), .Y(n10210) );
  AOI21XL U20122 ( .A0(n10209), .A1(n10245), .B0(n10210), .Y(n10211) );
  INVXL U20123 ( .A(n10213), .Y(n10215) );
  INVXL U20124 ( .A(n10219), .Y(n10221) );
  NAND2XL U20125 ( .A(n10234), .B(n10229), .Y(n10236) );
  OAI21XL U20126 ( .A0(n10231), .A1(n10195), .B0(n10230), .Y(n10232) );
  INVXL U20127 ( .A(n10237), .Y(n10239) );
  INVXL U20128 ( .A(n10240), .Y(n10242) );
  INVXL U20129 ( .A(n10209), .Y(n10241) );
  OAI21XL U20130 ( .A0(n10267), .A1(n10266), .B0(n10269), .Y(n10248) );
  OAI21XL U20131 ( .A0(M2_U4_U1_enc_tree_2__4__16_), .A1(
        M2_U3_U1_enc_tree_2__4__16_), .B0(n10248), .Y(n10255) );
  INVXL U20132 ( .A(n10279), .Y(n10281) );
  INVXL U20133 ( .A(n10283), .Y(n10285) );
  OAI22XL U20134 ( .A0(n10296), .A1(n10324), .B0(n10326), .B1(n10295), .Y(
        n10343) );
  XNOR2XL U20135 ( .A(n10494), .B(n10335), .Y(n10331) );
  OAI22XL U20136 ( .A0(n10517), .A1(n10299), .B0(n10533), .B1(n10331), .Y(
        n10348) );
  XNOR2X1 U20137 ( .A(n4808), .B(n10539), .Y(n10323) );
  OAI22XL U20138 ( .A0(n9504), .A1(n10301), .B0(n10496), .B1(n10323), .Y(
        n10346) );
  XNOR2XL U20139 ( .A(n10339), .B(M2_mult_x_15_n1668), .Y(n10327) );
  OAI22XL U20140 ( .A0(n10368), .A1(n10308), .B0(n10369), .B1(n10327), .Y(
        n10357) );
  XNOR2XL U20141 ( .A(M2_mult_x_15_n43), .B(n10515), .Y(n10328) );
  OAI22XL U20142 ( .A0(n4570), .A1(n10309), .B0(n10403), .B1(n10328), .Y(
        n10356) );
  CMPR32X1 U20143 ( .A(n10312), .B(n10311), .C(n10310), .CO(n10355), .S(n10314) );
  CMPR32X1 U20144 ( .A(n10315), .B(n10314), .C(n10313), .CO(n10431), .S(n10292) );
  INVXL U20145 ( .A(n10465), .Y(n10321) );
  NAND2X1 U20146 ( .A(n10320), .B(n10319), .Y(n10463) );
  XNOR2X1 U20147 ( .A(M2_a_17_), .B(n10538), .Y(n10334) );
  OAI22XL U20148 ( .A0(n9504), .A1(n10323), .B0(n10496), .B1(n10334), .Y(
        n10354) );
  OAI2BB1XL U20149 ( .A0N(n10326), .A1N(n10325), .B0(n10324), .Y(n10353) );
  OAI22XL U20150 ( .A0(n10368), .A1(n10327), .B0(n10369), .B1(n10339), .Y(
        n10352) );
  OAI22X1 U20151 ( .A0(n10541), .A1(n10330), .B0(n3174), .B1(n10336), .Y(
        n10350) );
  XNOR2X1 U20152 ( .A(n10494), .B(n10514), .Y(n10332) );
  OAI22XL U20153 ( .A0(n10532), .A1(n10331), .B0(n10533), .B1(n10332), .Y(
        n10349) );
  XNOR2X1 U20154 ( .A(n10494), .B(n10539), .Y(n10366) );
  OAI22XL U20155 ( .A0(n10517), .A1(n10332), .B0(n10533), .B1(n10366), .Y(
        n10372) );
  XNOR2XL U20156 ( .A(M2_mult_x_15_n43), .B(M2_mult_x_15_n1668), .Y(n10367) );
  XNOR2XL U20157 ( .A(n4808), .B(n10515), .Y(n10361) );
  OAI22XL U20158 ( .A0(n9504), .A1(n10334), .B0(n10496), .B1(n10361), .Y(
        n10370) );
  OAI22XL U20159 ( .A0(n10660), .A1(n10387), .B0(n3178), .B1(n10386), .Y(
        n10340) );
  OAI22XL U20160 ( .A0(n10368), .A1(n10339), .B0(n10369), .B1(n10338), .Y(
        n10363) );
  CMPR32X1 U20161 ( .A(n10351), .B(n10350), .C(n10349), .CO(n10411), .S(n10418) );
  CMPR32X1 U20162 ( .A(n10354), .B(n10353), .C(n10352), .CO(n10412), .S(n10417) );
  CMPR32X1 U20163 ( .A(n10357), .B(n10356), .C(n10355), .CO(n10416), .S(n10432) );
  XNOR2X1 U20164 ( .A(n4808), .B(M2_mult_x_15_n1669), .Y(n10381) );
  OAI22XL U20165 ( .A0(n9504), .A1(n10361), .B0(n10496), .B1(n10381), .Y(
        n10384) );
  OAI22XL U20166 ( .A0(n10660), .A1(n10337), .B0(n3178), .B1(M2_b_15_), .Y(
        n10385) );
  CMPR32X1 U20167 ( .A(n10372), .B(n10371), .C(n10370), .CO(n10373), .S(n10410) );
  XNOR2XL U20168 ( .A(n10494), .B(n10515), .Y(n10401) );
  OAI22XL U20169 ( .A0(n10532), .A1(n10380), .B0(n10533), .B1(n10401), .Y(
        n10399) );
  CMPR32X1 U20170 ( .A(n10384), .B(n10383), .C(n10382), .CO(n10408), .S(n10377) );
  CMPR32X1 U20171 ( .A(n10387), .B(n10386), .C(n10385), .CO(n10397), .S(n10382) );
  OAI22XL U20172 ( .A0(n10660), .A1(M2_b_15_), .B0(n3178), .B1(n10335), .Y(
        n10406) );
  CMPR32X1 U20173 ( .A(n10400), .B(n10399), .C(n10398), .CO(n10462), .S(n10409) );
  XNOR2XL U20174 ( .A(n10494), .B(M2_mult_x_15_n1669), .Y(n10457) );
  OAI22XL U20175 ( .A0(n10532), .A1(n10401), .B0(n10533), .B1(n10457), .Y(
        n10456) );
  OAI22XL U20176 ( .A0(n9504), .A1(n10404), .B0(n10496), .B1(n4808), .Y(n10452) );
  OAI22XL U20177 ( .A0(n10660), .A1(n10335), .B0(n10659), .B1(n10514), .Y(
        n10459) );
  CMPR32X1 U20178 ( .A(n6140), .B(n10406), .C(n10405), .CO(n10450), .S(n10396)
         );
  CMPR32X1 U20179 ( .A(n10409), .B(n10408), .C(n10407), .CO(n10447), .S(n10392) );
  CMPR32X1 U20180 ( .A(n10412), .B(n10411), .C(n10410), .CO(n10427), .S(n10442) );
  CMPR32X1 U20181 ( .A(n10415), .B(n10414), .C(n10413), .CO(n10423), .S(n10436) );
  CMPR32X1 U20182 ( .A(n10421), .B(n10420), .C(n10419), .CO(n10434), .S(n10439) );
  CMPR32X1 U20183 ( .A(n10424), .B(n10423), .C(n10422), .CO(n10426), .S(n10440) );
  CMPR32X1 U20184 ( .A(n10433), .B(n10432), .C(n10431), .CO(n10445), .S(n10437) );
  CMPR32X1 U20185 ( .A(n10449), .B(n10448), .C(n10447), .CO(n10482), .S(n10475) );
  CMPR32X1 U20186 ( .A(n10452), .B(n10451), .C(n10450), .CO(n10487), .S(n10460) );
  CMPR32X1 U20187 ( .A(n10456), .B(n10455), .C(n10454), .CO(n10498), .S(n10461) );
  OAI22XL U20188 ( .A0(n10517), .A1(n10457), .B0(n10533), .B1(n10495), .Y(
        n10490) );
  CMPR32X1 U20189 ( .A(n10337), .B(M2_b_15_), .C(n10459), .CO(n10488), .S(
        n10451) );
  CMPR32X1 U20190 ( .A(n10462), .B(n10461), .C(n10460), .CO(n10485), .S(n10448) );
  NOR2X1 U20191 ( .A(n10647), .B(n10521), .Y(n10639) );
  INVXL U20192 ( .A(n10639), .Y(n10484) );
  NAND2XL U20193 ( .A(n10469), .B(n10468), .Y(n10610) );
  INVXL U20194 ( .A(n10610), .Y(n10470) );
  NAND2XL U20195 ( .A(n10472), .B(n10471), .Y(n10607) );
  NAND2XL U20196 ( .A(n10476), .B(n10475), .Y(n10624) );
  OAI21XL U20197 ( .A0(n10623), .A1(n10630), .B0(n10624), .Y(n10477) );
  CMPR32X1 U20198 ( .A(n10487), .B(n10486), .C(n10485), .CO(n10502), .S(n10481) );
  CMPR32X1 U20199 ( .A(n10490), .B(n10489), .C(n10488), .CO(n10508), .S(n10497) );
  CMPR32X1 U20200 ( .A(n10499), .B(n10498), .C(n10497), .CO(n10506), .S(n10486) );
  CMPR32X1 U20201 ( .A(n10508), .B(n10507), .C(n10506), .CO(n10553), .S(n10501) );
  CMPR32X1 U20202 ( .A(n10511), .B(n10510), .C(n10509), .CO(n10524), .S(n10518) );
  XNOR2XL U20203 ( .A(n25885), .B(M2_mult_x_15_n1668), .Y(n10531) );
  CMPR32X1 U20204 ( .A(n10335), .B(n10514), .C(n10513), .CO(n10529), .S(n10520) );
  CMPR32X1 U20205 ( .A(n10520), .B(n10519), .C(n10518), .CO(n10522), .S(n10507) );
  NOR2X1 U20206 ( .A(n10553), .B(n10552), .Y(n10644) );
  INVX1 U20207 ( .A(n10644), .Y(n10555) );
  CMPR32X1 U20208 ( .A(n10527), .B(n10526), .C(n10525), .CO(n10536), .S(n10528) );
  CMPR32X1 U20209 ( .A(n10530), .B(n10529), .C(n10528), .CO(n10535), .S(n10523) );
  CMPR32X1 U20210 ( .A(n10536), .B(n10535), .C(n10534), .CO(n10560), .S(n10557) );
  CMPR32X1 U20211 ( .A(n10539), .B(n10538), .C(n10537), .CO(n10547), .S(n10542) );
  CMPR32X1 U20212 ( .A(n10544), .B(n10543), .C(n10542), .CO(n10545), .S(n10534) );
  CMPR32X1 U20213 ( .A(n10547), .B(n10546), .C(n10545), .CO(n10564), .S(n10559) );
  CMPR32X1 U20214 ( .A(n10516), .B(n10550), .C(n10549), .CO(n10567), .S(n10546) );
  NAND2XL U20215 ( .A(n10634), .B(n10646), .Y(n10566) );
  INVXL U20216 ( .A(n10645), .Y(n10554) );
  OAI21XL U20217 ( .A0(n10582), .A1(n10600), .B0(n10583), .Y(n10561) );
  AOI21XL U20218 ( .A0(n10635), .A1(n10646), .B0(n10651), .Y(n10565) );
  OAI21X1 U20219 ( .A0(n5237), .A1(n10566), .B0(n10565), .Y(n10573) );
  CMPR32X1 U20220 ( .A(n10569), .B(n10568), .C(n10567), .CO(n10572), .S(n10563) );
  CMPR32X1 U20221 ( .A(n10515), .B(M2_mult_x_15_n1669), .C(n10570), .CO(n10657), .S(n10568) );
  NOR2X1 U20222 ( .A(n10647), .B(n10578), .Y(n10596) );
  INVXL U20223 ( .A(n10576), .Y(n10577) );
  INVXL U20224 ( .A(n10586), .Y(n10587) );
  AOI21X1 U20225 ( .A0(n10635), .A1(n10588), .B0(n10587), .Y(n10589) );
  INVXL U20226 ( .A(n10596), .Y(n10599) );
  OAI21X2 U20227 ( .A0(n5237), .A1(n10599), .B0(n10598), .Y(n10602) );
  INVXL U20228 ( .A(n10603), .Y(n10613) );
  NAND2XL U20229 ( .A(n10612), .B(n10613), .Y(n10606) );
  INVXL U20230 ( .A(n10604), .Y(n10616) );
  AOI21XL U20231 ( .A0(n10503), .A1(n10613), .B0(n10616), .Y(n10605) );
  NAND2XL U20232 ( .A(n10612), .B(n10505), .Y(n10609) );
  NAND2XL U20233 ( .A(n10626), .B(n10631), .Y(n10622) );
  AOI21X1 U20234 ( .A0(n10616), .A1(n4619), .B0(n10615), .Y(n10617) );
  INVXL U20235 ( .A(n10630), .Y(n10620) );
  INVXL U20236 ( .A(n10626), .Y(n10629) );
  NAND2X1 U20237 ( .A(n10631), .B(n10630), .Y(n10632) );
  INVXL U20238 ( .A(n10635), .Y(n10636) );
  NAND2XL U20239 ( .A(n10639), .B(n10641), .Y(n10643) );
  OR2X2 U20240 ( .A(n10647), .B(n10653), .Y(n10655) );
  CMPR32X1 U20241 ( .A(n3177), .B(n10658), .C(n10657), .CO(n10663), .S(n10571)
         );
  CLKINVX3 U20242 ( .A(n20993), .Y(n23722) );
  OAI21XL U20243 ( .A0(n10708), .A1(n10707), .B0(n10706), .Y(n10710) );
  INVXL U20244 ( .A(n23492), .Y(n10714) );
  NOR2XL U20245 ( .A(n10714), .B(n10713), .Y(n10715) );
  BUFX3 U20246 ( .A(n10719), .Y(n25807) );
  AND2X2 U20247 ( .A(n2982), .B(n23967), .Y(n25723) );
  AOI21XL U20248 ( .A0(n10722), .A1(n23862), .B0(n10721), .Y(n10723) );
  NOR2XL U20249 ( .A(n20279), .B(n20275), .Y(n10740) );
  NOR2XL U20250 ( .A(M6_mult_x_15_n717), .B(M6_mult_x_15_n721), .Y(n10897) );
  OAI21X1 U20251 ( .A0(n11057), .A1(n25895), .B0(n10746), .Y(n11168) );
  OAI21XL U20252 ( .A0(n11057), .A1(n25896), .B0(n10747), .Y(n11163) );
  OAI21X1 U20253 ( .A0(n11057), .A1(n26226), .B0(n10750), .Y(n11166) );
  CLKINVX3 U20254 ( .A(n22989), .Y(n22987) );
  INVX1 U20255 ( .A(n11216), .Y(n22490) );
  NOR2X4 U20256 ( .A(n10760), .B(n10759), .Y(n23023) );
  AND3X2 U20257 ( .A(n10760), .B(n10759), .C(n10758), .Y(n23021) );
  OAI21XL U20258 ( .A0(n22978), .A1(n23025), .B0(n10761), .Y(n10762) );
  INVX1 U20259 ( .A(n11209), .Y(n22614) );
  XOR2XL U20260 ( .A(n10762), .B(n3054), .Y(n23218) );
  INVXL U20261 ( .A(n11131), .Y(n10763) );
  NAND2X1 U20262 ( .A(n10763), .B(n10771), .Y(n22985) );
  OAI2BB2XL U20263 ( .B0(n22886), .B1(n3225), .A0N(n22987), .A1N(n22887), .Y(
        n10764) );
  INVXL U20264 ( .A(n10764), .Y(n10765) );
  OAI21XL U20265 ( .A0(n22985), .A1(n23025), .B0(n10765), .Y(n10766) );
  OAI21XL U20266 ( .A0(n23025), .A1(n22989), .B0(n10767), .Y(n10768) );
  NOR2X1 U20267 ( .A(n11163), .B(n11165), .Y(n11139) );
  OAI22X1 U20268 ( .A0(n11057), .A1(n26217), .B0(n9107), .B1(n25951), .Y(
        n11162) );
  NAND2XL U20269 ( .A(n10852), .B(n10850), .Y(n10776) );
  NOR2X4 U20270 ( .A(n10785), .B(n10784), .Y(n22932) );
  AND3X2 U20271 ( .A(n10785), .B(n10784), .C(n10783), .Y(n22931) );
  AOI222XL U20272 ( .A0(n22932), .A1(n10775), .B0(n22904), .B1(n10769), .C0(
        n22931), .C1(n23002), .Y(n10786) );
  OAI21XL U20273 ( .A0(n22993), .A1(n22912), .B0(n10786), .Y(n10787) );
  XOR2XL U20274 ( .A(n10787), .B(n3053), .Y(n10884) );
  OAI21XL U20275 ( .A0(n10872), .A1(n11047), .B0(n11049), .Y(n10792) );
  AOI222XL U20276 ( .A0(n22953), .A1(n10789), .B0(n10797), .B1(n3220), .C0(
        n22952), .C1(n26496), .Y(n10800) );
  OAI21XL U20277 ( .A0(n23148), .A1(n22834), .B0(n10800), .Y(n10801) );
  NOR2XL U20278 ( .A(M6_mult_x_15_n722), .B(n10894), .Y(n10802) );
  NOR2XL U20279 ( .A(n10897), .B(n10802), .Y(n10900) );
  AOI222XL U20280 ( .A0(n22953), .A1(n10775), .B0(n10797), .B1(n10769), .C0(
        n22952), .C1(n23002), .Y(n10803) );
  OAI21XL U20281 ( .A0(n22993), .A1(n22834), .B0(n10803), .Y(n10804) );
  XOR2XL U20282 ( .A(n10804), .B(n3221), .Y(n10838) );
  AOI222XL U20283 ( .A0(n22932), .A1(n10749), .B0(n22904), .B1(n3116), .C0(
        n22931), .C1(n22987), .Y(n10805) );
  OAI21XL U20284 ( .A0(n22978), .A1(n22912), .B0(n10805), .Y(n10806) );
  XOR2XL U20285 ( .A(n10806), .B(n3053), .Y(n10849) );
  INVXL U20286 ( .A(n10807), .Y(n10808) );
  OAI21XL U20287 ( .A0(n22985), .A1(n22912), .B0(n10808), .Y(n10809) );
  XOR2XL U20288 ( .A(n10809), .B(n3053), .Y(n10820) );
  OAI21XL U20289 ( .A0(n22912), .A1(n22989), .B0(n4709), .Y(n10810) );
  XOR2XL U20290 ( .A(n10810), .B(n11216), .Y(n10829) );
  NOR2XL U20291 ( .A(n10838), .B(n10837), .Y(n10841) );
  OAI21XL U20292 ( .A0(n11139), .A1(n10824), .B0(n10822), .Y(n10816) );
  NAND2XL U20293 ( .A(n10814), .B(n10813), .Y(n10815) );
  AOI222XL U20294 ( .A0(n22953), .A1(n10769), .B0(n10797), .B1(n23002), .C0(
        n22952), .C1(n10749), .Y(n10817) );
  OAI21XL U20295 ( .A0(n22998), .A1(n22834), .B0(n10817), .Y(n10818) );
  XOR2XL U20296 ( .A(n10818), .B(n3221), .Y(n10836) );
  CMPR22X1 U20297 ( .A(n10820), .B(n10819), .CO(n10848), .S(n10835) );
  NOR2XL U20298 ( .A(n10836), .B(n10835), .Y(n10821) );
  NOR2XL U20299 ( .A(n10841), .B(n10821), .Y(n10844) );
  AOI222XL U20300 ( .A0(n22953), .A1(n23002), .B0(n10797), .B1(n10749), .C0(
        n22952), .C1(n3116), .Y(n10826) );
  OAI21XL U20301 ( .A0(n23006), .A1(n22834), .B0(n10826), .Y(n10827) );
  XOR2XL U20302 ( .A(n10827), .B(n3221), .Y(n10831) );
  INVXL U20303 ( .A(n10831), .Y(n10834) );
  NOR3XL U20304 ( .A(n22987), .B(n10749), .C(n3116), .Y(n10828) );
  NAND2XL U20305 ( .A(n10828), .B(n3221), .Y(n10833) );
  CMPR22X1 U20306 ( .A(n3053), .B(n10829), .CO(n10819), .S(n10830) );
  NAND2XL U20307 ( .A(n10831), .B(n10830), .Y(n10832) );
  OAI21XL U20308 ( .A0(n10834), .A1(n10833), .B0(n10832), .Y(n10843) );
  NAND2XL U20309 ( .A(n10836), .B(n10835), .Y(n10840) );
  NAND2XL U20310 ( .A(n10838), .B(n10837), .Y(n10839) );
  OAI21XL U20311 ( .A0(n10841), .A1(n10840), .B0(n10839), .Y(n10842) );
  AOI21XL U20312 ( .A0(n10844), .A1(n10843), .B0(n10842), .Y(n10865) );
  CMPR22X1 U20313 ( .A(n3054), .B(n10845), .CO(n10866), .S(n10877) );
  AOI222XL U20314 ( .A0(n22932), .A1(n23002), .B0(n22904), .B1(n10749), .C0(
        n22931), .C1(n3116), .Y(n10846) );
  OAI21XL U20315 ( .A0(n23006), .A1(n22912), .B0(n10846), .Y(n10847) );
  XOR2XL U20316 ( .A(n10847), .B(n3053), .Y(n10876) );
  ADDHXL U20317 ( .A(n10849), .B(n10848), .CO(n10875), .S(n10837) );
  AOI222XL U20318 ( .A0(n22953), .A1(n26496), .B0(n10797), .B1(n10775), .C0(
        n22952), .C1(n10769), .Y(n10859) );
  OAI21XL U20319 ( .A0(n22924), .A1(n22834), .B0(n10859), .Y(n10860) );
  XOR2XL U20320 ( .A(n10860), .B(n3221), .Y(n10861) );
  NOR2XL U20321 ( .A(n10862), .B(n10861), .Y(n10864) );
  NAND2XL U20322 ( .A(n10862), .B(n10861), .Y(n10863) );
  OAI21XL U20323 ( .A0(n10865), .A1(n10864), .B0(n10863), .Y(n10882) );
  CMPR22X1 U20324 ( .A(n10867), .B(n10866), .CO(n23217), .S(n10888) );
  AOI222XL U20325 ( .A0(n22932), .A1(n10769), .B0(n22904), .B1(n23002), .C0(
        n22931), .C1(n10749), .Y(n10868) );
  OAI21XL U20326 ( .A0(n22998), .A1(n22912), .B0(n10868), .Y(n10869) );
  XOR2XL U20327 ( .A(n10869), .B(n3053), .Y(n10887) );
  AOI222XL U20328 ( .A0(n22953), .A1(n3220), .B0(n10797), .B1(n22867), .C0(
        n22952), .C1(n10775), .Y(n10873) );
  OAI21XL U20329 ( .A0(n22869), .A1(n22834), .B0(n10873), .Y(n10874) );
  XOR2XL U20330 ( .A(n10874), .B(n3221), .Y(n10886) );
  CMPR32X1 U20331 ( .A(n10877), .B(n10876), .C(n10875), .CO(n10878), .S(n10862) );
  OR2XL U20332 ( .A(n10879), .B(n10878), .Y(n10881) );
  AND2XL U20333 ( .A(n10879), .B(n10878), .Y(n10880) );
  AOI21XL U20334 ( .A0(n10882), .A1(n10881), .B0(n10880), .Y(n10893) );
  CMPR32X1 U20335 ( .A(n10885), .B(n10884), .C(n10883), .CO(n10894), .S(n10890) );
  CMPR32X1 U20336 ( .A(n10888), .B(n10887), .C(n10886), .CO(n10889), .S(n10879) );
  NOR2XL U20337 ( .A(n10890), .B(n10889), .Y(n10892) );
  NAND2XL U20338 ( .A(n10890), .B(n10889), .Y(n10891) );
  OAI21XL U20339 ( .A0(n10893), .A1(n10892), .B0(n10891), .Y(n10899) );
  NAND2XL U20340 ( .A(M6_mult_x_15_n722), .B(n10894), .Y(n10896) );
  NAND2XL U20341 ( .A(M6_mult_x_15_n717), .B(M6_mult_x_15_n721), .Y(n10895) );
  OAI21XL U20342 ( .A0(n10897), .A1(n10896), .B0(n10895), .Y(n10898) );
  NOR2XL U20343 ( .A(M6_mult_x_15_n712), .B(M6_mult_x_15_n716), .Y(n10902) );
  NAND2XL U20344 ( .A(M6_mult_x_15_n712), .B(M6_mult_x_15_n716), .Y(n10901) );
  OAI21XL U20345 ( .A0(n10903), .A1(n10902), .B0(n10901), .Y(n10910) );
  NOR2XL U20346 ( .A(M6_mult_x_15_n698), .B(M6_mult_x_15_n704), .Y(n10907) );
  NOR2XL U20347 ( .A(M6_mult_x_15_n705), .B(M6_mult_x_15_n711), .Y(n10904) );
  NOR2XL U20348 ( .A(n10907), .B(n10904), .Y(n10909) );
  NAND2XL U20349 ( .A(M6_mult_x_15_n705), .B(M6_mult_x_15_n711), .Y(n10906) );
  NAND2XL U20350 ( .A(M6_mult_x_15_n698), .B(M6_mult_x_15_n704), .Y(n10905) );
  OAI21XL U20351 ( .A0(n10907), .A1(n10906), .B0(n10905), .Y(n10908) );
  AOI21XL U20352 ( .A0(n10910), .A1(n10909), .B0(n10908), .Y(n10917) );
  OR2XL U20353 ( .A(M6_mult_x_15_n683), .B(M6_mult_x_15_n690), .Y(n10914) );
  OR2XL U20354 ( .A(M6_mult_x_15_n691), .B(M6_mult_x_15_n697), .Y(n10911) );
  NAND2XL U20355 ( .A(n10914), .B(n10911), .Y(n10916) );
  AND2XL U20356 ( .A(M6_mult_x_15_n691), .B(M6_mult_x_15_n697), .Y(n10913) );
  AND2XL U20357 ( .A(M6_mult_x_15_n683), .B(M6_mult_x_15_n690), .Y(n10912) );
  AOI21XL U20358 ( .A0(n10914), .A1(n10913), .B0(n10912), .Y(n10915) );
  OAI21XL U20359 ( .A0(n10917), .A1(n10916), .B0(n10915), .Y(n10924) );
  NOR2XL U20360 ( .A(M6_mult_x_15_n675), .B(M6_mult_x_15_n682), .Y(n10918) );
  NOR2XL U20361 ( .A(n10921), .B(n10918), .Y(n10923) );
  NAND2XL U20362 ( .A(M6_mult_x_15_n675), .B(M6_mult_x_15_n682), .Y(n10920) );
  NAND2XL U20363 ( .A(M6_mult_x_15_n667), .B(M6_mult_x_15_n674), .Y(n10919) );
  OAI21XL U20364 ( .A0(n10921), .A1(n10920), .B0(n10919), .Y(n10922) );
  OAI21XL U20365 ( .A0(n10930), .A1(n10929), .B0(n10928), .Y(n10935) );
  OAI21XL U20366 ( .A0(n10933), .A1(n10932), .B0(n10931), .Y(n10934) );
  OAI21XL U20367 ( .A0(n11126), .A1(n11276), .B0(n11127), .Y(n11107) );
  OAI21XL U20368 ( .A0(n11109), .A1(n11120), .B0(n11110), .Y(n10937) );
  OAI21XL U20369 ( .A0(n10940), .A1(n11106), .B0(n10939), .Y(n10983) );
  OAI21XL U20370 ( .A0(n11101), .A1(n11115), .B0(n11102), .Y(n11039) );
  OAI21XL U20371 ( .A0(n11340), .A1(n11336), .B0(n11341), .Y(n10941) );
  OAI21XL U20372 ( .A0(n11031), .A1(n11345), .B0(n11032), .Y(n10987) );
  OAI21XL U20373 ( .A0(n10992), .A1(n11096), .B0(n10993), .Y(n10943) );
  OAI21XL U20374 ( .A0(n10984), .A1(n10946), .B0(n10945), .Y(n10947) );
  OAI21XL U20375 ( .A0(n11357), .A1(n11354), .B0(n11358), .Y(n11023) );
  OAI21XL U20376 ( .A0(n10979), .A1(n10973), .B0(n10974), .Y(n11018) );
  OAI21XL U20377 ( .A0(n10961), .A1(n10959), .B0(n11008), .Y(n10958) );
  OAI21XL U20378 ( .A0(n10963), .A1(n10962), .B0(n10968), .Y(n10967) );
  OAI21XL U20379 ( .A0(n10972), .A1(n10978), .B0(n10979), .Y(n10977) );
  OAI21XL U20380 ( .A0(n11118), .A1(n10985), .B0(n10984), .Y(n11030) );
  OAI21XL U20381 ( .A0(n11348), .A1(n10989), .B0(n10988), .Y(n11099) );
  OAI21XL U20382 ( .A0(n10998), .A1(n10997), .B0(n11350), .Y(n11002) );
  OAI21XL U20383 ( .A0(n11015), .A1(n11014), .B0(n11013), .Y(n11016) );
  AOI21XL U20384 ( .A0(n11018), .A1(n11017), .B0(n11016), .Y(n11019) );
  OAI21XL U20385 ( .A0(n11021), .A1(n11020), .B0(n11019), .Y(n11022) );
  AOI21XL U20386 ( .A0(n11372), .A1(n11026), .B0(n11025), .Y(n11045) );
  NAND2XL U20387 ( .A(n11362), .B(n11364), .Y(n11027) );
  OAI21XL U20388 ( .A0(n11118), .A1(n11041), .B0(n11040), .Y(n11339) );
  OAI21XL U20389 ( .A0(n11045), .A1(n11044), .B0(n11364), .Y(n11095) );
  OAI21XL U20390 ( .A0(n11056), .A1(n11055), .B0(n11054), .Y(n21085) );
  OAI22X1 U20391 ( .A0(n23193), .A1(n26224), .B0(n9107), .B1(n25943), .Y(
        n11149) );
  INVX1 U20392 ( .A(n11149), .Y(n22549) );
  OAI22X1 U20393 ( .A0(n11057), .A1(n25991), .B0(n9107), .B1(n25891), .Y(
        n11157) );
  NOR2X1 U20394 ( .A(n11155), .B(n11157), .Y(n22642) );
  INVX1 U20395 ( .A(n11157), .Y(n22636) );
  OAI21XL U20396 ( .A0(n22584), .A1(n11067), .B0(n11066), .Y(n11068) );
  OAI21XL U20397 ( .A0(n22504), .A1(n11079), .B0(n11078), .Y(n21067) );
  INVX1 U20398 ( .A(n11169), .Y(n21056) );
  NAND2BX2 U20399 ( .AN(n21057), .B(n21056), .Y(n23154) );
  AND3X2 U20400 ( .A(n21057), .B(n11090), .C(n21056), .Y(n23150) );
  OAI21XL U20401 ( .A0(n11082), .A1(n11089), .B0(n11091), .Y(n11092) );
  NAND2XL U20402 ( .A(n11367), .B(n11365), .Y(n11094) );
  OAI21XL U20403 ( .A0(n11118), .A1(n11114), .B0(n11115), .Y(n11105) );
  OAI21XL U20404 ( .A0(n11123), .A1(n11119), .B0(n11120), .Y(n11113) );
  OR4XL U20405 ( .A(n23022), .B(n11151), .C(n11147), .D(n11149), .Y(n11237) );
  AOI21XL U20406 ( .A0(n22553), .A1(n22500), .B0(n11237), .Y(n11132) );
  NOR4X1 U20407 ( .A(n11160), .B(n11162), .C(n22867), .D(n11159), .Y(n11239)
         );
  NAND2XL U20408 ( .A(n22642), .B(n22605), .Y(n11238) );
  NAND2XL U20409 ( .A(n11131), .B(n11139), .Y(n11240) );
  AOI221XL U20410 ( .A0(n11132), .A1(n11239), .B0(n11238), .B1(n11239), .C0(
        n11240), .Y(n11268) );
  OAI21XL U20411 ( .A0(n23089), .A1(n11133), .B0(n22500), .Y(n11134) );
  AOI211XL U20412 ( .A0(n22553), .A1(n11134), .B0(n11147), .C0(n11149), .Y(
        n11135) );
  OAI31XL U20413 ( .A0(n23022), .A1(n11151), .A2(n11135), .B0(n22605), .Y(
        n11136) );
  AOI211XL U20414 ( .A0(n22642), .A1(n11136), .B0(n22867), .C0(n11159), .Y(
        n11137) );
  OR3XL U20415 ( .A(n11160), .B(n11162), .C(n11137), .Y(n11138) );
  INVXL U20416 ( .A(n11210), .Y(n11170) );
  AOI21XL U20417 ( .A0(n11170), .A1(n11169), .B0(n22713), .Y(n11176) );
  INVXL U20418 ( .A(n22491), .Y(n11175) );
  OAI21XL U20419 ( .A0(n11176), .A1(n22492), .B0(n11175), .Y(n11181) );
  AOI21XL U20420 ( .A0(n11181), .A1(n22698), .B0(n21059), .Y(n11186) );
  INVXL U20421 ( .A(n21062), .Y(n11191) );
  OAI21XL U20422 ( .A0(n11192), .A1(n21063), .B0(n11191), .Y(n11197) );
  INVX1 U20423 ( .A(n21089), .Y(n22967) );
  AOI21XL U20424 ( .A0(n11197), .A1(n22967), .B0(n21078), .Y(n11200) );
  OAI21XL U20425 ( .A0(n11200), .A1(n21079), .B0(n22614), .Y(n11202) );
  INVXL U20426 ( .A(n11214), .Y(n11201) );
  AOI21XL U20427 ( .A0(n11202), .A1(n11201), .B0(n11213), .Y(n11204) );
  INVXL U20428 ( .A(n11217), .Y(n11203) );
  OAI21XL U20429 ( .A0(n11204), .A1(n11216), .B0(n11203), .Y(n11206) );
  INVXL U20430 ( .A(n11219), .Y(n11205) );
  AOI21XL U20431 ( .A0(n11206), .A1(n11205), .B0(n11220), .Y(n11208) );
  OAI21XL U20432 ( .A0(n11208), .A1(n11221), .B0(n11207), .Y(n11453) );
  NOR2XL U20433 ( .A(n21079), .B(n11209), .Y(n11229) );
  NOR2XL U20434 ( .A(n21062), .B(n21063), .Y(n11225) );
  NOR2XL U20435 ( .A(n22716), .B(n21059), .Y(n11227) );
  NOR2XL U20436 ( .A(n22492), .B(n22491), .Y(n11228) );
  OAI21XL U20437 ( .A0(n11210), .A1(n22713), .B0(n11228), .Y(n11211) );
  NOR2XL U20438 ( .A(n21058), .B(n22990), .Y(n11226) );
  OAI2BB1XL U20439 ( .A0N(n11227), .A1N(n11211), .B0(n11226), .Y(n11212) );
  NOR2XL U20440 ( .A(n21078), .B(n21089), .Y(n11230) );
  OAI2BB1XL U20441 ( .A0N(n11225), .A1N(n11212), .B0(n11230), .Y(n11215) );
  NOR2XL U20442 ( .A(n11214), .B(n11213), .Y(n11232) );
  OAI2BB1XL U20443 ( .A0N(n11229), .A1N(n11215), .B0(n11232), .Y(n11218) );
  NOR2XL U20444 ( .A(n11217), .B(n11216), .Y(n11231) );
  NAND2XL U20445 ( .A(n11218), .B(n11231), .Y(n11224) );
  NOR2XL U20446 ( .A(n11220), .B(n11219), .Y(n11235) );
  NOR2XL U20447 ( .A(n11222), .B(n11221), .Y(n11234) );
  INVXL U20448 ( .A(n11234), .Y(n11223) );
  AOI21XL U20449 ( .A0(n11224), .A1(n11235), .B0(n11223), .Y(n11269) );
  NAND2XL U20450 ( .A(n11226), .B(n11225), .Y(n11241) );
  AOI21XL U20451 ( .A0(n11228), .A1(n11227), .B0(n11241), .Y(n11233) );
  NAND2XL U20452 ( .A(n11230), .B(n11229), .Y(n11242) );
  NAND2XL U20453 ( .A(n11232), .B(n11231), .Y(n11244) );
  AOI2BB1XL U20454 ( .A0N(n11233), .A1N(n11242), .B0(n11244), .Y(n11236) );
  NAND2XL U20455 ( .A(n11235), .B(n11234), .Y(n11243) );
  NOR2XL U20456 ( .A(n11236), .B(n11243), .Y(n11266) );
  NOR2XL U20457 ( .A(n11238), .B(n11237), .Y(n11252) );
  NAND2BXL U20458 ( .AN(n11240), .B(n11239), .Y(n11251) );
  NOR2XL U20459 ( .A(n11252), .B(n11251), .Y(n11247) );
  OR2XL U20460 ( .A(n11242), .B(n11241), .Y(n11248) );
  NOR2XL U20461 ( .A(n11244), .B(n11243), .Y(n11250) );
  NAND2XL U20462 ( .A(n11248), .B(n11250), .Y(n11246) );
  INVXL U20463 ( .A(n11246), .Y(n11245) );
  AND2XL U20464 ( .A(n11247), .B(n11245), .Y(n11254) );
  NAND2BXL U20465 ( .AN(n11247), .B(n11246), .Y(n11255) );
  OAI21XL U20466 ( .A0(n11257), .A1(n11254), .B0(n11255), .Y(n11259) );
  INVXL U20467 ( .A(n11248), .Y(n11249) );
  NAND2XL U20468 ( .A(n11250), .B(n11249), .Y(n11264) );
  INVXL U20469 ( .A(n11264), .Y(n11253) );
  AOI21XL U20470 ( .A0(n11275), .A1(n11253), .B0(n11265), .Y(n11263) );
  NOR2BXL U20471 ( .AN(n11255), .B(n11254), .Y(n11256) );
  INVXL U20472 ( .A(n11258), .Y(n11262) );
  NAND2BXL U20473 ( .AN(n11265), .B(n11264), .Y(n11274) );
  CMPR32X1 U20474 ( .A(n11268), .B(n11267), .C(n11266), .CO(n11257), .S(n11272) );
  CMPR32X1 U20475 ( .A(n11270), .B(n11450), .C(n11269), .CO(n11267), .S(n11271) );
  OAI21XL U20476 ( .A0(n11275), .A1(n11274), .B0(n11273), .Y(n11451) );
  NAND2XL U20477 ( .A(n11311), .B(y10[30]), .Y(n11281) );
  NAND2XL U20478 ( .A(n9106), .B(y11[30]), .Y(n11280) );
  NAND2XL U20479 ( .A(n11311), .B(y10[29]), .Y(n11283) );
  NAND2XL U20480 ( .A(n9106), .B(y11[29]), .Y(n11282) );
  MXI2X1 U20481 ( .A(w2[61]), .B(w2[93]), .S0(valid[0]), .Y(n11437) );
  NAND2XL U20482 ( .A(w2[56]), .B(n23973), .Y(n11285) );
  NAND2XL U20483 ( .A(w2[88]), .B(valid[0]), .Y(n11284) );
  NAND2XL U20484 ( .A(w2[55]), .B(n23973), .Y(n11287) );
  NAND2XL U20485 ( .A(w2[87]), .B(valid[0]), .Y(n11286) );
  MXI2X1 U20486 ( .A(w2[57]), .B(w2[89]), .S0(valid[0]), .Y(n11440) );
  NAND2XL U20487 ( .A(w2[58]), .B(n23973), .Y(n11289) );
  NAND2XL U20488 ( .A(w2[90]), .B(valid[0]), .Y(n11288) );
  MXI2X1 U20489 ( .A(w2[59]), .B(w2[91]), .S0(valid[0]), .Y(n11435) );
  NAND2XL U20490 ( .A(w2[60]), .B(n23973), .Y(n11291) );
  NAND2XL U20491 ( .A(w2[92]), .B(valid[0]), .Y(n11290) );
  NAND2XL U20492 ( .A(n11311), .B(y10[28]), .Y(n11293) );
  NAND2XL U20493 ( .A(n9106), .B(y11[28]), .Y(n11292) );
  OAI21XL U20494 ( .A0(n11298), .A1(n11434), .B0(n11294), .Y(n11295) );
  NAND2XL U20495 ( .A(n11311), .B(y10[27]), .Y(n11297) );
  NAND2XL U20496 ( .A(n9106), .B(y11[27]), .Y(n11296) );
  NAND2XL U20497 ( .A(n11311), .B(y10[26]), .Y(n11300) );
  NAND2XL U20498 ( .A(n9106), .B(y11[26]), .Y(n11299) );
  OAI21XL U20499 ( .A0(n11305), .A1(n11439), .B0(n11301), .Y(n11302) );
  NAND2XL U20500 ( .A(n11311), .B(y10[25]), .Y(n11304) );
  NAND2XL U20501 ( .A(n9106), .B(y11[25]), .Y(n11303) );
  NAND2XL U20502 ( .A(n11311), .B(y10[24]), .Y(n11307) );
  NAND2XL U20503 ( .A(n9106), .B(y11[24]), .Y(n11306) );
  NAND2XL U20504 ( .A(n11307), .B(n11306), .Y(n11428) );
  INVXL U20505 ( .A(n11308), .Y(n11310) );
  NOR2XL U20506 ( .A(n11309), .B(n11326), .Y(n11442) );
  NOR2XL U20507 ( .A(n11310), .B(n11442), .Y(n11325) );
  NAND2XL U20508 ( .A(n11311), .B(y10[23]), .Y(n11313) );
  NAND2XL U20509 ( .A(n9106), .B(y11[23]), .Y(n11312) );
  NAND2XL U20510 ( .A(n11313), .B(n11312), .Y(n11413) );
  INVXL U20511 ( .A(n11413), .Y(n11429) );
  NOR2XL U20512 ( .A(n11429), .B(n11326), .Y(n11324) );
  NAND2XL U20513 ( .A(w2[62]), .B(n23973), .Y(n11315) );
  NAND2XL U20514 ( .A(w2[94]), .B(valid[0]), .Y(n11314) );
  CMPR32X1 U20515 ( .A(n11418), .B(n11317), .C(n11316), .CO(n11400), .S(n25835) );
  CMPR32X1 U20516 ( .A(n11421), .B(n11319), .C(n11318), .CO(n11316), .S(n24443) );
  CMPR32X1 U20517 ( .A(n11427), .B(n11321), .C(n11320), .CO(n11328), .S(n25716) );
  CMPR32X1 U20518 ( .A(n11426), .B(n11323), .C(n11322), .CO(n11320), .S(n23786) );
  CMPR32X1 U20519 ( .A(n11428), .B(n11325), .C(n11324), .CO(n11322), .S(n25704) );
  INVXL U20520 ( .A(n11326), .Y(n11327) );
  XOR2XL U20521 ( .A(n11413), .B(n11327), .Y(n25701) );
  NOR4XL U20522 ( .A(n25716), .B(n23786), .C(n25704), .D(n25701), .Y(n11330)
         );
  CMPR32X1 U20523 ( .A(n11420), .B(n11329), .C(n11328), .CO(n11318), .S(n25072) );
  INVXL U20524 ( .A(n25072), .Y(n11405) );
  NAND4BXL U20525 ( .AN(n11349), .B(n11459), .C(n11473), .D(n11468), .Y(n11380) );
  AOI21XL U20526 ( .A0(n11372), .A1(n11356), .B0(n11355), .Y(n11361) );
  OAI21XL U20527 ( .A0(n11371), .A1(n11370), .B0(n11369), .Y(n11390) );
  AOI21XL U20528 ( .A0(n11372), .A1(n11386), .B0(n11390), .Y(n11379) );
  INVX1 U20529 ( .A(n11082), .Y(n22913) );
  OAI21XL U20530 ( .A0(n22913), .A1(n23154), .B0(n11373), .Y(n11374) );
  CMPR32X1 U20531 ( .A(n11395), .B(M6_mult_x_15_n433), .C(n11375), .CO(n11376), 
        .S(n11093) );
  NAND2XL U20532 ( .A(n11389), .B(n11387), .Y(n11378) );
  NAND4BXL U20533 ( .AN(n11380), .B(n20289), .C(n23599), .D(n20721), .Y(n11381) );
  OAI21XL U20534 ( .A0(n11393), .A1(n11392), .B0(n11391), .Y(n11398) );
  CMPR32X1 U20535 ( .A(n11071), .B(n11395), .C(n11394), .CO(n11396), .S(n11377) );
  CMPR32X1 U20536 ( .A(n11419), .B(n11400), .C(n11401), .CO(n11402), .S(n23678) );
  INVXL U20537 ( .A(n25835), .Y(n11406) );
  INVXL U20538 ( .A(n23786), .Y(n11404) );
  NAND2XL U20539 ( .A(n25704), .B(n25701), .Y(n23785) );
  NAND4XL U20540 ( .A(n25072), .B(n25716), .C(n25704), .D(n23786), .Y(n11408)
         );
  NAND4XL U20541 ( .A(n11418), .B(n11419), .C(n11420), .D(n11421), .Y(n11417)
         );
  NAND4XL U20542 ( .A(n11426), .B(n11427), .C(n11428), .D(n11413), .Y(n11416)
         );
  NAND2XL U20543 ( .A(n11414), .B(n11433), .Y(n11415) );
  OAI21XL U20544 ( .A0(n11417), .A1(n11416), .B0(n11415), .Y(n25245) );
  INVXL U20545 ( .A(n11418), .Y(n11425) );
  INVXL U20546 ( .A(n11419), .Y(n11424) );
  INVXL U20547 ( .A(n11420), .Y(n11423) );
  INVXL U20548 ( .A(n11421), .Y(n11422) );
  NAND4XL U20549 ( .A(n11425), .B(n11424), .C(n11423), .D(n11422), .Y(n11446)
         );
  INVXL U20550 ( .A(n11426), .Y(n11432) );
  INVXL U20551 ( .A(n11427), .Y(n11431) );
  INVXL U20552 ( .A(n11428), .Y(n11430) );
  NAND4XL U20553 ( .A(n11432), .B(n11431), .C(n11430), .D(n11429), .Y(n11445)
         );
  INVXL U20554 ( .A(n11433), .Y(n11438) );
  INVXL U20555 ( .A(n11434), .Y(n11436) );
  NAND4XL U20556 ( .A(n11438), .B(n11437), .C(n11436), .D(n11435), .Y(n11444)
         );
  INVXL U20557 ( .A(n11439), .Y(n11441) );
  NAND3XL U20558 ( .A(n11442), .B(n11441), .C(n11440), .Y(n11443) );
  CLKINVX3 U20559 ( .A(n20717), .Y(n23949) );
  INVXL U20560 ( .A(n11449), .Y(n11452) );
  OAI21XL U20561 ( .A0(n19064), .A1(n20959), .B0(n19065), .Y(n11464) );
  CLKINVX3 U20562 ( .A(n20728), .Y(n23947) );
  AOI22XL U20563 ( .A0(n23949), .A1(n23919), .B0(n23947), .B1(n23886), .Y(
        n11476) );
  OAI22X1 U20564 ( .A0(n6211), .A1(n15942), .B0(n25899), .B1(n25813), .Y(
        n11491) );
  BUFX3 U20565 ( .A(n11491), .Y(M3_mult_x_15_b_14_) );
  OAI21X2 U20566 ( .A0(n25813), .A1(n26248), .B0(n11492), .Y(M3_a_9_) );
  OAI22X1 U20567 ( .A0(n26025), .A1(n4860), .B0(n25898), .B1(n25796), .Y(
        n11496) );
  OAI222X1 U20568 ( .A0(n25909), .A1(n4860), .B0(n26258), .B1(n25813), .C0(
        n26009), .C1(n15940), .Y(M3_a_0_) );
  OAI222X1 U20569 ( .A0(n6187), .A1(n15942), .B0(n25910), .B1(n25813), .C0(
        n15940), .C1(n23989), .Y(n11497) );
  AOI21XL U20570 ( .A0(n14417), .A1(y11[7]), .B0(n25145), .Y(n11500) );
  OAI21XL U20571 ( .A0(n25243), .A1(n25897), .B0(n11500), .Y(M1_a_7_) );
  CLKINVX3 U20572 ( .A(n13720), .Y(n25860) );
  AOI21XL U20573 ( .A0(n14417), .A1(y11[6]), .B0(n25144), .Y(n11502) );
  OAI21XL U20574 ( .A0(n25243), .A1(n25906), .B0(n11502), .Y(M1_a_6_) );
  AOI21XL U20575 ( .A0(n14417), .A1(y11[1]), .B0(n25139), .Y(n11503) );
  OAI21XL U20576 ( .A0(n25243), .A1(n25898), .B0(n11503), .Y(M1_a_1_) );
  AOI21XL U20577 ( .A0(n14417), .A1(y11[0]), .B0(n24266), .Y(n11506) );
  OAI21X1 U20578 ( .A0(n25243), .A1(n25909), .B0(n11506), .Y(M1_a_0_) );
  AOI21XL U20579 ( .A0(n14417), .A1(y11[5]), .B0(n25143), .Y(n11507) );
  OAI21XL U20580 ( .A0(n25243), .A1(n25902), .B0(n11507), .Y(M1_a_5_) );
  AOI22XL U20581 ( .A0(n4566), .A1(learning_rate[4]), .B0(in_valid_d), .B1(
        w1[132]), .Y(n11509) );
  AOI21XL U20582 ( .A0(n14417), .A1(y11[4]), .B0(n25142), .Y(n11510) );
  NAND2X1 U20583 ( .A(n11512), .B(n11511), .Y(M1_b_6_) );
  AOI21XL U20584 ( .A0(n14417), .A1(y11[2]), .B0(n25140), .Y(n11513) );
  AOI22XL U20585 ( .A0(n4566), .A1(learning_rate[0]), .B0(in_valid_d), .B1(
        w1[128]), .Y(n11515) );
  NAND2X1 U20586 ( .A(n11515), .B(n11514), .Y(M1_b_0_) );
  AOI21XL U20587 ( .A0(n14417), .A1(y11[9]), .B0(n25147), .Y(n11516) );
  AOI21XL U20588 ( .A0(n14417), .A1(y11[8]), .B0(n25146), .Y(n11517) );
  AOI21XL U20589 ( .A0(n14417), .A1(y11[3]), .B0(n25141), .Y(n11518) );
  AOI21XL U20590 ( .A0(n14417), .A1(y11[10]), .B0(n25148), .Y(n11519) );
  OAI21XL U20591 ( .A0(n25243), .A1(n25905), .B0(n11519), .Y(M1_a_10_) );
  AOI22XL U20592 ( .A0(n11536), .A1(learning_rate[10]), .B0(in_valid_d), .B1(
        w1[138]), .Y(n11521) );
  AOI21XL U20593 ( .A0(n14417), .A1(y11[11]), .B0(n25149), .Y(n11523) );
  AOI21XL U20594 ( .A0(n14417), .A1(y11[12]), .B0(n25150), .Y(n11524) );
  AOI21XL U20595 ( .A0(n14417), .A1(y11[13]), .B0(n25151), .Y(n11525) );
  AOI21XL U20596 ( .A0(n14417), .A1(y11[14]), .B0(n25152), .Y(n11526) );
  NAND2X1 U20597 ( .A(in_valid_d), .B(w1[143]), .Y(n11528) );
  INVX8 U20598 ( .A(n14197), .Y(n25862) );
  NAND2X1 U20599 ( .A(n11530), .B(n11529), .Y(M1_b_14_) );
  AOI21XL U20600 ( .A0(n14417), .A1(y11[15]), .B0(n25153), .Y(n11532) );
  AOI21XL U20601 ( .A0(n14417), .A1(y11[16]), .B0(n25154), .Y(n11535) );
  AOI22XL U20602 ( .A0(n11536), .A1(learning_rate[18]), .B0(in_valid_d), .B1(
        w1[146]), .Y(n11538) );
  AOI21XL U20603 ( .A0(n14417), .A1(y11[17]), .B0(n25155), .Y(n11539) );
  NAND2X1 U20604 ( .A(n3123), .B(w1[147]), .Y(n11542) );
  OAI21XL U20605 ( .A0(n25243), .A1(n25914), .B0(n3557), .Y(M1_a_19_) );
  AOI21XL U20606 ( .A0(n14417), .A1(y11[21]), .B0(n25158), .Y(n11545) );
  OAI21XL U20607 ( .A0(n25243), .A1(n25913), .B0(n11545), .Y(M1_a_21_) );
  AOI21XL U20608 ( .A0(n14417), .A1(y11[22]), .B0(n24024), .Y(n11548) );
  OAI21XL U20609 ( .A0(n25243), .A1(n25915), .B0(n11548), .Y(M1_a_22_) );
  OAI21XL U20610 ( .A0(n26046), .A1(n15940), .B0(n11552), .Y(n11554) );
  OAI21XL U20611 ( .A0(n26037), .A1(n17167), .B0(n11555), .Y(n11557) );
  NOR2X1 U20612 ( .A(n11557), .B(n11556), .Y(n13004) );
  OAI21XL U20613 ( .A0(n26036), .A1(n17167), .B0(n11558), .Y(n11560) );
  OAI21XL U20614 ( .A0(n26043), .A1(n15940), .B0(n11564), .Y(n11566) );
  OAI21XL U20615 ( .A0(n26301), .A1(n15940), .B0(n11570), .Y(n11572) );
  XOR2X1 U20616 ( .A(n13004), .B(n13005), .Y(n11610) );
  NAND3X2 U20617 ( .A(n11602), .B(n11601), .C(n11600), .Y(n18780) );
  CMPR32X1 U20618 ( .A(n18770), .B(n11606), .C(n11605), .CO(n11603), .S(n25789) );
  CMPR32X1 U20619 ( .A(n18773), .B(n11608), .C(n11607), .CO(n11615), .S(n25184) );
  CMPR32X1 U20620 ( .A(n18779), .B(n11610), .C(n11609), .CO(n11611), .S(n24087) );
  CMPR32X1 U20621 ( .A(n18776), .B(n11612), .C(n11611), .CO(n11607), .S(n24336) );
  CMPR22X1 U20622 ( .A(n13004), .B(n18780), .CO(n11609), .S(n25804) );
  CMPR32X1 U20623 ( .A(n18783), .B(n11614), .C(n11613), .CO(n11605), .S(n24376) );
  NAND4BXL U20624 ( .AN(n25789), .B(n11619), .C(n11618), .D(n11617), .Y(n11620) );
  NOR3X1 U20625 ( .A(n24040), .B(n25791), .C(n11620), .Y(n12940) );
  NAND2BX1 U20626 ( .AN(n24040), .B(n11623), .Y(n24046) );
  XNOR2X1 U20627 ( .A(n25884), .B(n3190), .Y(n11641) );
  OAI22X1 U20628 ( .A0(n12357), .A1(n11652), .B0(n12284), .B1(n12282), .Y(
        n11668) );
  OAI22XL U20629 ( .A0(n12152), .A1(n11653), .B0(n3185), .B1(n11635), .Y(
        n11667) );
  XNOR2X1 U20630 ( .A(n12233), .B(M5_b_18_), .Y(n11648) );
  XNOR2X1 U20631 ( .A(n12233), .B(M3_mult_x_15_b_19_), .Y(n11637) );
  NAND2X4 U20632 ( .A(n11627), .B(n12746), .Y(n12715) );
  XNOR2X1 U20633 ( .A(n12732), .B(n3049), .Y(n11663) );
  XNOR2X1 U20634 ( .A(n12732), .B(n3197), .Y(n11629) );
  INVX4 U20635 ( .A(M3_mult_x_15_a_17_), .Y(n12696) );
  XNOR2X1 U20636 ( .A(M3_mult_x_15_a_17_), .B(M3_mult_x_15_b_9_), .Y(n11639)
         );
  OAI22XL U20637 ( .A0(n12717), .A1(n11649), .B0(n12718), .B1(n11639), .Y(
        n11665) );
  XNOR2X1 U20638 ( .A(n12519), .B(n12560), .Y(n11687) );
  OAI22XL U20639 ( .A0(n12635), .A1(n11687), .B0(n12633), .B1(n11642), .Y(
        n11632) );
  INVX4 U20640 ( .A(M3_mult_x_15_n61), .Y(n12751) );
  XNOR2X1 U20641 ( .A(n12758), .B(n3108), .Y(n11689) );
  XNOR2X1 U20642 ( .A(n12758), .B(n3049), .Y(n11643) );
  OAI22X1 U20643 ( .A0(n12759), .A1(n11689), .B0(n12760), .B1(n11643), .Y(
        n11631) );
  XNOR2X1 U20644 ( .A(n3204), .B(M5_b_18_), .Y(n11654) );
  XNOR2X1 U20645 ( .A(M3_mult_x_15_a_17_), .B(n16884), .Y(n11638) );
  OAI22XL U20646 ( .A0(n12717), .A1(n11638), .B0(n12718), .B1(n11762), .Y(
        n11772) );
  XNOR2X1 U20647 ( .A(n25884), .B(n12561), .Y(n11640) );
  XNOR2XL U20648 ( .A(n12265), .B(n3202), .Y(n11634) );
  OAI22XL U20649 ( .A0(n12352), .A1(n11636), .B0(n12222), .B1(n11763), .Y(
        n11759) );
  XOR2X1 U20650 ( .A(M3_a_10_), .B(M3_a_11_), .Y(n11633) );
  INVX8 U20651 ( .A(n12522), .Y(n12594) );
  XNOR2X1 U20652 ( .A(n12594), .B(n3198), .Y(n11647) );
  XNOR2X1 U20653 ( .A(n12594), .B(n3021), .Y(n11695) );
  OAI22XL U20654 ( .A0(n12597), .A1(n11647), .B0(n12523), .B1(n11695), .Y(
        n11708) );
  OAI22X1 U20655 ( .A0(n12357), .A1(n12282), .B0(n3183), .B1(n12285), .Y(
        n11707) );
  OAI22XL U20656 ( .A0(n12152), .A1(n11635), .B0(n3185), .B1(n11634), .Y(
        n11706) );
  OAI22X1 U20657 ( .A0(n12352), .A1(n11637), .B0(n12222), .B1(n11636), .Y(
        n11705) );
  OAI22X2 U20658 ( .A0(n12717), .A1(n11639), .B0(n12718), .B1(n11638), .Y(
        n11704) );
  OAI22XL U20659 ( .A0(n12618), .A1(n11641), .B0(n12119), .B1(n11640), .Y(
        n11703) );
  OAI22X1 U20660 ( .A0(n12759), .A1(n11643), .B0(n12760), .B1(n11782), .Y(
        n11779) );
  OAI2BB1XL U20661 ( .A0N(n12284), .A1N(n12025), .B0(n12282), .Y(n11778) );
  XNOR2X1 U20662 ( .A(n3204), .B(n3198), .Y(n11673) );
  XNOR2X1 U20663 ( .A(n3204), .B(n3021), .Y(n11644) );
  OAI22X1 U20664 ( .A0(n12535), .A1(n3110), .B0(n12995), .B1(M3_mult_x_15_b_1_), .Y(n11675) );
  XNOR2X1 U20665 ( .A(n3204), .B(n3201), .Y(n11655) );
  OAI22XL U20666 ( .A0(n12597), .A1(n11650), .B0(n12523), .B1(n11647), .Y(
        n11656) );
  NAND2X1 U20667 ( .A(n2980), .B(n4775), .Y(n12293) );
  XNOR2X1 U20668 ( .A(n12732), .B(n3108), .Y(n11664) );
  OAI22XL U20669 ( .A0(n12715), .A1(n11744), .B0(n12525), .B1(n11664), .Y(
        n11729) );
  XNOR2X1 U20670 ( .A(n25884), .B(M3_mult_x_15_b_9_), .Y(n11723) );
  OAI22X1 U20671 ( .A0(n12618), .A1(n11723), .B0(n12119), .B1(n11651), .Y(
        n11685) );
  XNOR2XL U20672 ( .A(n12265), .B(M3_mult_x_15_b_19_), .Y(n11672) );
  OAI22XL U20673 ( .A0(n12152), .A1(n11672), .B0(n3185), .B1(n11653), .Y(
        n11683) );
  OAI22XL U20674 ( .A0(n12598), .A1(n11655), .B0(n12342), .B1(n11654), .Y(
        n11700) );
  CMPR32X1 U20675 ( .A(n11658), .B(n11657), .C(n11656), .CO(n11698), .S(n11659) );
  OAI22XL U20676 ( .A0(n12635), .A1(n11670), .B0(n12513), .B1(n11688), .Y(
        n11679) );
  OAI22X1 U20677 ( .A0(n12759), .A1(n11662), .B0(n12760), .B1(n11690), .Y(
        n11678) );
  OAI22XL U20678 ( .A0(n12715), .A1(n11664), .B0(n12525), .B1(n11663), .Y(
        n11677) );
  OAI22X1 U20679 ( .A0(n12357), .A1(n11793), .B0(n3183), .B1(n11671), .Y(
        n11800) );
  XNOR2XL U20680 ( .A(n12265), .B(M5_b_18_), .Y(n11795) );
  OAI22XL U20681 ( .A0(n12152), .A1(n11795), .B0(n3185), .B1(n11672), .Y(
        n11799) );
  XNOR2XL U20682 ( .A(n3204), .B(n12701), .Y(n11747) );
  OAI22XL U20683 ( .A0(n12598), .A1(n11747), .B0(n12342), .B1(n11673), .Y(
        n11733) );
  XNOR2X1 U20684 ( .A(M3_a_11_), .B(n3201), .Y(n11764) );
  OAI22XL U20685 ( .A0(n12597), .A1(n11695), .B0(n12523), .B1(n11764), .Y(
        n11777) );
  OAI22XL U20686 ( .A0(n12535), .A1(n11499), .B0(n12995), .B1(n3108), .Y(
        n11765) );
  CMPR32X1 U20687 ( .A(n11700), .B(n11699), .C(n11698), .CO(n11770), .S(n11694) );
  ADDFHX1 U20688 ( .A(n11702), .B(n11701), .CI(n11691), .CO(n11714), .S(n11709) );
  ADDFHX1 U20689 ( .A(n11708), .B(n11707), .CI(n11706), .CO(n11758), .S(n11712) );
  OAI22XL U20690 ( .A0(n12352), .A1(n11746), .B0(n12222), .B1(n11721), .Y(
        n11798) );
  XNOR2X1 U20691 ( .A(n12716), .B(n3108), .Y(n11829) );
  XNOR2X1 U20692 ( .A(n3204), .B(n12560), .Y(n11831) );
  OAI22XL U20693 ( .A0(n12598), .A1(n11831), .B0(n12342), .B1(n11747), .Y(
        n11808) );
  OAI22XL U20694 ( .A0(n12576), .A1(n12751), .B0(n11749), .B1(n11748), .Y(
        n11817) );
  XNOR2X1 U20695 ( .A(n12519), .B(M3_mult_x_15_b_9_), .Y(n11792) );
  XNOR2X1 U20696 ( .A(n12282), .B(M5_b_18_), .Y(n11851) );
  XNOR2X1 U20697 ( .A(n12265), .B(n3201), .Y(n11796) );
  OAI22XL U20698 ( .A0(n12152), .A1(n11847), .B0(n3185), .B1(n11796), .Y(
        n11853) );
  XNOR2X1 U20699 ( .A(n12716), .B(n12561), .Y(n11877) );
  XNOR2X1 U20700 ( .A(n12233), .B(n3202), .Y(n11892) );
  OAI22X2 U20701 ( .A0(n12352), .A1(n11763), .B0(n12222), .B1(n11892), .Y(
        n11884) );
  XOR3X2 U20702 ( .A(n11883), .B(n11884), .C(n11887), .Y(n11897) );
  XNOR2X1 U20703 ( .A(n12594), .B(M5_b_18_), .Y(n11876) );
  OAI22XL U20704 ( .A0(n12597), .A1(n11764), .B0(n12523), .B1(n11876), .Y(
        n11895) );
  CMPR32X1 U20705 ( .A(M3_mult_x_15_b_1_), .B(n12279), .C(n11765), .CO(n11893), 
        .S(n11775) );
  ADDFHX4 U20706 ( .A(n11768), .B(n11767), .CI(n11766), .CO(n11900), .S(n11786) );
  ADDFHX1 U20707 ( .A(n11780), .B(n11779), .CI(n11778), .CO(n11888), .S(n11756) );
  ADDFHX1 U20708 ( .A(n11801), .B(n11800), .CI(n11799), .CO(n11742), .S(n11820) );
  CMPR32X1 U20709 ( .A(n11810), .B(n11809), .C(n11808), .CO(n11837), .S(n12446) );
  XNOR2X1 U20710 ( .A(n12594), .B(n16884), .Y(n11842) );
  XNOR2X1 U20711 ( .A(n12758), .B(n3110), .Y(n11813) );
  OAI22XL U20712 ( .A0(n12618), .A1(n11844), .B0(n12119), .B1(n11816), .Y(
        n12450) );
  XNOR2X1 U20713 ( .A(n2980), .B(M3_mult_x_15_b_19_), .Y(n11848) );
  OAI22X1 U20714 ( .A0(n12340), .A1(n11848), .B0(n11819), .B1(n12338), .Y(
        n11999) );
  XNOR2X1 U20715 ( .A(n12594), .B(M3_mult_x_15_b_9_), .Y(n12001) );
  OAI22XL U20716 ( .A0(n12597), .A1(n12001), .B0(n12595), .B1(n11842), .Y(
        n12048) );
  XNOR2X1 U20717 ( .A(M3_mult_x_15_a_17_), .B(n12279), .Y(n12004) );
  XNOR2X1 U20718 ( .A(n25884), .B(n3108), .Y(n12026) );
  OAI22XL U20719 ( .A0(n12618), .A1(n12026), .B0(n12119), .B1(n11844), .Y(
        n12046) );
  XNOR2X1 U20720 ( .A(n12265), .B(n3198), .Y(n11992) );
  OAI22XL U20721 ( .A0(n12152), .A1(n11992), .B0(n3185), .B1(n11847), .Y(
        n12051) );
  XNOR2XL U20722 ( .A(n12233), .B(n12560), .Y(n11994) );
  XNOR2X1 U20723 ( .A(n2980), .B(M5_b_18_), .Y(n11997) );
  OAI22XL U20724 ( .A0(n12340), .A1(n11997), .B0(n11848), .B1(n4775), .Y(
        n11996) );
  OAI22XL U20725 ( .A0(n12715), .A1(n12731), .B0(n12525), .B1(n11849), .Y(
        n11995) );
  XNOR2X1 U20726 ( .A(n3204), .B(n3190), .Y(n12021) );
  OAI22XL U20727 ( .A0(n12598), .A1(n12021), .B0(n12342), .B1(n11850), .Y(
        n12008) );
  XNOR2X1 U20728 ( .A(n12282), .B(n3201), .Y(n12023) );
  OAI22X1 U20729 ( .A0(n12357), .A1(n12023), .B0(n12284), .B1(n11851), .Y(
        n12007) );
  OAI22XL U20730 ( .A0(n12635), .A1(n11993), .B0(n12513), .B1(n11852), .Y(
        n12006) );
  ADDFHX2 U20731 ( .A(n11860), .B(n11859), .CI(n11858), .CO(n11865), .S(n12472) );
  ADDFHX4 U20732 ( .A(n11863), .B(n11862), .CI(n11861), .CO(n12500), .S(n12499) );
  CMPR32X1 U20733 ( .A(n11869), .B(n11868), .C(n11867), .CO(n11904), .S(n11901) );
  OAI22XL U20734 ( .A0(n12597), .A1(n11876), .B0(n12523), .B1(n11926), .Y(
        n11925) );
  OAI22XL U20735 ( .A0(n12635), .A1(n11878), .B0(n12633), .B1(n11915), .Y(
        n11923) );
  OAI22XL U20736 ( .A0(n12715), .A1(n11880), .B0(n12525), .B1(n11918), .Y(
        n11921) );
  OAI22XL U20737 ( .A0(n12535), .A1(n3049), .B0(n12995), .B1(n3197), .Y(n11927) );
  INVXL U20738 ( .A(n11883), .Y(n11882) );
  NAND2BXL U20739 ( .AN(n11884), .B(n11882), .Y(n11886) );
  ADDFHX1 U20740 ( .A(n11889), .B(n11888), .CI(n4658), .CO(n11933), .S(n11873)
         );
  OAI2BB1XL U20741 ( .A0N(n3185), .A1N(n12152), .B0(n12265), .Y(n11911) );
  CMPR32X1 U20742 ( .A(n11895), .B(n11894), .C(n11893), .CO(n11908), .S(n11896) );
  CMPR32X1 U20743 ( .A(n11907), .B(n11906), .C(n11905), .CO(n11936), .S(n11928) );
  OAI22XL U20744 ( .A0(n12635), .A1(n11915), .B0(n12633), .B1(n11951), .Y(
        n11943) );
  INVX4 U20745 ( .A(n12696), .Y(n12716) );
  XNOR2X1 U20746 ( .A(n12716), .B(n12701), .Y(n11946) );
  OAI22X1 U20747 ( .A0(n12578), .A1(n11916), .B0(n12718), .B1(n11946), .Y(
        n11956) );
  CMPR32X1 U20748 ( .A(n11925), .B(n11924), .C(n11923), .CO(n11941), .S(n11930) );
  OAI22XL U20749 ( .A0(n12597), .A1(n11926), .B0(n12523), .B1(n11950), .Y(
        n11949) );
  CMPR32X1 U20750 ( .A(n11499), .B(n3108), .C(n11927), .CO(n11948), .S(n11907)
         );
  OAI22XL U20751 ( .A0(n12352), .A1(n12233), .B0(n12222), .B1(n11486), .Y(
        n11952) );
  CMPR32X1 U20752 ( .A(n11930), .B(n11929), .C(n11928), .CO(n11938), .S(n11920) );
  ADDFHX1 U20753 ( .A(n11933), .B(n11931), .CI(n11932), .CO(n11937), .S(n11919) );
  CMPR32X1 U20754 ( .A(n11936), .B(n11935), .C(n11934), .CO(n11967), .S(n11964) );
  ADDFHX1 U20755 ( .A(n11939), .B(n11938), .CI(n11937), .CO(n11966), .S(n11962) );
  XNOR2X1 U20756 ( .A(n12758), .B(n3190), .Y(n11984) );
  XNOR2X1 U20757 ( .A(n12716), .B(n3198), .Y(n11978) );
  OAI22XL U20758 ( .A0(n12578), .A1(n11946), .B0(n12718), .B1(n11978), .Y(
        n11976) );
  CMPR32X1 U20759 ( .A(n11949), .B(n11948), .C(n11947), .CO(n11974), .S(n11940) );
  XNOR2X1 U20760 ( .A(n12594), .B(n12803), .Y(n11979) );
  OAI22XL U20761 ( .A0(n12597), .A1(n11950), .B0(n12523), .B1(n11979), .Y(
        n11983) );
  OAI22XL U20762 ( .A0(n12535), .A1(M3_mult_x_15_n1682), .B0(n12995), .B1(
        M3_mult_x_15_b_9_), .Y(n11986) );
  OAI22XL U20763 ( .A0(n12598), .A1(n11958), .B0(n12342), .B1(n3204), .Y(
        n11988) );
  ADDFHX1 U20764 ( .A(n11967), .B(n11966), .CI(n11965), .CO(n12512), .S(n12510) );
  XNOR2X1 U20765 ( .A(n12716), .B(n3021), .Y(n12593) );
  OAI22XL U20766 ( .A0(n11979), .A1(n12597), .B0(n12523), .B1(n12596), .Y(
        n12629) );
  OAI22XL U20767 ( .A0(n12635), .A1(n11980), .B0(n12633), .B1(n12634), .Y(
        n12628) );
  XNOR2XL U20768 ( .A(n25884), .B(M5_b_18_), .Y(n12617) );
  XNOR2XL U20769 ( .A(n12758), .B(n12561), .Y(n12637) );
  OAI22XL U20770 ( .A0(n12598), .A1(n3204), .B0(n12342), .B1(n12225), .Y(
        n12620) );
  XNOR2XL U20771 ( .A(n12265), .B(n12701), .Y(n12011) );
  OAI22XL U20772 ( .A0(n12152), .A1(n12011), .B0(n3185), .B1(n11992), .Y(
        n12054) );
  XNOR2X1 U20773 ( .A(n12519), .B(n3049), .Y(n12013) );
  OAI22XL U20774 ( .A0(n12352), .A1(n12033), .B0(n12222), .B1(n11994), .Y(
        n12052) );
  ADDHXL U20775 ( .A(n11996), .B(n11995), .CO(n12049), .S(n12060) );
  NOR2BX1 U20776 ( .AN(n3110), .B(n12525), .Y(n12039) );
  XNOR2X1 U20777 ( .A(n2980), .B(n3201), .Y(n12031) );
  OAI22X1 U20778 ( .A0(n12340), .A1(n12031), .B0(n11997), .B1(n12338), .Y(
        n12038) );
  OAI22XL U20779 ( .A0(n12357), .A1(n12010), .B0(n12284), .B1(n12024), .Y(
        n12014) );
  OAI22X1 U20780 ( .A0(n12717), .A1(n12005), .B0(n12718), .B1(n12004), .Y(
        n12020) );
  XNOR2X1 U20781 ( .A(n12594), .B(n3049), .Y(n12072) );
  XNOR2X1 U20782 ( .A(n12265), .B(n12561), .Y(n12071) );
  OAI22XL U20783 ( .A0(n12152), .A1(n12071), .B0(n3185), .B1(n12012), .Y(
        n12067) );
  OAI22XL U20784 ( .A0(n12598), .A1(n12030), .B0(n12342), .B1(n12022), .Y(
        n12019) );
  OAI22X1 U20785 ( .A0(n12152), .A1(n12012), .B0(n3185), .B1(n12011), .Y(
        n12018) );
  XNOR2X1 U20786 ( .A(n12519), .B(n3108), .Y(n12029) );
  OAI22XL U20787 ( .A0(n12635), .A1(n12029), .B0(n12513), .B1(n12013), .Y(
        n12017) );
  ADDFHX1 U20788 ( .A(n12016), .B(n12015), .CI(n12014), .CO(n12058), .S(n12080) );
  ADDFHX1 U20789 ( .A(n12019), .B(n12018), .CI(n12017), .CO(n12042), .S(n12081) );
  OAI22XL U20790 ( .A0(n12598), .A1(n12022), .B0(n12342), .B1(n12021), .Y(
        n12045) );
  OAI22X1 U20791 ( .A0(n12025), .A1(n12024), .B0(n12284), .B1(n12023), .Y(
        n12044) );
  OAI22XL U20792 ( .A0(n12618), .A1(n12027), .B0(n12119), .B1(n12026), .Y(
        n12043) );
  XNOR2X1 U20793 ( .A(M3_mult_x_15_a_17_), .B(n3110), .Y(n12028) );
  OAI22XL U20794 ( .A0(n12635), .A1(n12066), .B0(n12513), .B1(n12029), .Y(
        n12074) );
  XNOR2X1 U20795 ( .A(n12233), .B(n3190), .Y(n12034) );
  OAI22XL U20796 ( .A0(n12352), .A1(n12073), .B0(n12222), .B1(n12034), .Y(
        n12079) );
  OAI22X1 U20797 ( .A0(n12578), .A1(n12696), .B0(n12718), .B1(n12032), .Y(
        n12035) );
  CMPR32X1 U20798 ( .A(n12051), .B(n12050), .C(n12049), .CO(n12436), .S(n12454) );
  XNOR2X1 U20799 ( .A(n25884), .B(M3_mult_x_15_b_1_), .Y(n12100) );
  XNOR2X1 U20800 ( .A(n3204), .B(n3197), .Y(n12099) );
  XNOR2X1 U20801 ( .A(n12519), .B(n12279), .Y(n12102) );
  ADDFHX1 U20802 ( .A(n12069), .B(n12068), .CI(n12067), .CO(n12082), .S(n12103) );
  OAI22XL U20803 ( .A0(n12152), .A1(n12117), .B0(n3185), .B1(n12071), .Y(
        n12110) );
  OAI22XL U20804 ( .A0(n12352), .A1(n12106), .B0(n12222), .B1(n12073), .Y(
        n12108) );
  CMPR32X1 U20805 ( .A(n12079), .B(n12078), .C(n12077), .CO(n12090), .S(n12114) );
  ADDFHX1 U20806 ( .A(n12082), .B(n12081), .CI(n12080), .CO(n12085), .S(n12092) );
  XNOR2X1 U20807 ( .A(n2980), .B(n12701), .Y(n12120) );
  ADDFHX1 U20808 ( .A(n12098), .B(n12097), .CI(n12096), .CO(n12104), .S(n12123) );
  XNOR2XL U20809 ( .A(n3204), .B(n3049), .Y(n12125) );
  OAI22XL U20810 ( .A0(n12598), .A1(n12125), .B0(n12342), .B1(n12099), .Y(
        n12130) );
  XNOR2X1 U20811 ( .A(n25884), .B(n3110), .Y(n12101) );
  OAI22X1 U20812 ( .A0(n12618), .A1(n12101), .B0(n12119), .B1(n12100), .Y(
        n12129) );
  OAI22XL U20813 ( .A0(n12635), .A1(n12121), .B0(n12513), .B1(n12102), .Y(
        n12128) );
  XNOR2X1 U20814 ( .A(n12282), .B(n12561), .Y(n12127) );
  OAI22XL U20815 ( .A0(n12357), .A1(n12127), .B0(n12284), .B1(n12105), .Y(
        n12143) );
  XNOR2XL U20816 ( .A(n12594), .B(n11499), .Y(n12126) );
  XNOR2X1 U20817 ( .A(n12233), .B(n5430), .Y(n12131) );
  OAI22XL U20818 ( .A0(n12352), .A1(n12131), .B0(n12222), .B1(n12106), .Y(
        n12141) );
  ADDFHX1 U20819 ( .A(n12110), .B(n12109), .CI(n12108), .CO(n12116), .S(n12138) );
  OAI22XL U20820 ( .A0(n12635), .A1(n12163), .B0(n12513), .B1(n12121), .Y(
        n12147) );
  XNOR2X1 U20821 ( .A(n12594), .B(n12279), .Y(n12165) );
  OAI22XL U20822 ( .A0(n12357), .A1(n12150), .B0(n12284), .B1(n12127), .Y(
        n12153) );
  XNOR2X1 U20823 ( .A(n12265), .B(M3_mult_x_15_b_9_), .Y(n12151) );
  XNOR2X1 U20824 ( .A(n12233), .B(n3197), .Y(n12162) );
  XNOR2X1 U20825 ( .A(n2980), .B(n12561), .Y(n12170) );
  OAI22XL U20826 ( .A0(n12635), .A1(M3_U3_U1_or2_inv_0__18_), .B0(n12513), 
        .B1(n12132), .Y(n12169) );
  CMPR32X1 U20827 ( .A(n12137), .B(n12136), .C(n12135), .CO(n12423), .S(n12422) );
  ADDFHX1 U20828 ( .A(n12149), .B(n12148), .CI(n12147), .CO(n12144), .S(n12180) );
  XNOR2X1 U20829 ( .A(n12282), .B(n16884), .Y(n12173) );
  XNOR2X1 U20830 ( .A(n12265), .B(n5430), .Y(n12174) );
  OAI22XL U20831 ( .A0(n12152), .A1(n12174), .B0(n3185), .B1(n12151), .Y(
        n12184) );
  XNOR2X1 U20832 ( .A(n12233), .B(n3049), .Y(n12172) );
  XNOR2X1 U20833 ( .A(n12519), .B(n3110), .Y(n12164) );
  XNOR2X1 U20834 ( .A(n12594), .B(n12271), .Y(n12171) );
  OAI22XL U20835 ( .A0(n12597), .A1(n12171), .B0(n12595), .B1(n12165), .Y(
        n12181) );
  NOR2BX1 U20836 ( .AN(n3110), .B(n12513), .Y(n12190) );
  XNOR2X1 U20837 ( .A(n2980), .B(n3190), .Y(n12186) );
  OAI22X1 U20838 ( .A0(n12340), .A1(n12186), .B0(n12170), .B1(n12338), .Y(
        n12189) );
  XNOR2X1 U20839 ( .A(n12233), .B(n3108), .Y(n12200) );
  OAI22XL U20840 ( .A0(n12352), .A1(n12200), .B0(n12222), .B1(n12172), .Y(
        n12209) );
  XNOR2X1 U20841 ( .A(n12282), .B(M3_mult_x_15_b_9_), .Y(n12203) );
  OAI22X1 U20842 ( .A0(n12357), .A1(n12203), .B0(n12284), .B1(n12173), .Y(
        n12208) );
  XNOR2XL U20843 ( .A(n12265), .B(n3197), .Y(n12204) );
  OAI22XL U20844 ( .A0(n12152), .A1(n12204), .B0(n3185), .B1(n12174), .Y(
        n12207) );
  ADDFHX1 U20845 ( .A(n12180), .B(n12179), .CI(n12178), .CO(n12175), .S(n12196) );
  CMPR32X1 U20846 ( .A(n12183), .B(n12182), .C(n12181), .CO(n12193), .S(n12212) );
  ADDFHX1 U20847 ( .A(n12190), .B(n12189), .CI(n12188), .CO(n12198), .S(n12388) );
  NOR2X1 U20848 ( .A(n12411), .B(n12410), .Y(n12414) );
  OAI22XL U20849 ( .A0(n12352), .A1(n12350), .B0(n12222), .B1(n12200), .Y(
        n12360) );
  XNOR2X1 U20850 ( .A(n12594), .B(n3110), .Y(n12202) );
  OAI22XL U20851 ( .A0(n12597), .A1(n12202), .B0(n12595), .B1(n12201), .Y(
        n12359) );
  XNOR2X1 U20852 ( .A(n12282), .B(n5430), .Y(n12355) );
  OAI22XL U20853 ( .A0(n12357), .A1(n12355), .B0(n12284), .B1(n12203), .Y(
        n12358) );
  XNOR2X1 U20854 ( .A(n12265), .B(n3049), .Y(n12353) );
  OAI22XL U20855 ( .A0(n12152), .A1(n12353), .B0(n3185), .B1(n12204), .Y(
        n12335) );
  CMPR32X1 U20856 ( .A(n12212), .B(n12211), .C(n12210), .CO(n12195), .S(n12385) );
  NOR2XL U20857 ( .A(n12409), .B(n12408), .Y(n12213) );
  NOR2XL U20858 ( .A(n12414), .B(n12213), .Y(n12218) );
  XNOR2X1 U20859 ( .A(n12233), .B(n12279), .Y(n12351) );
  OAI22XL U20860 ( .A0(n12352), .A1(n12228), .B0(n12222), .B1(n12351), .Y(
        n12346) );
  XNOR2X1 U20861 ( .A(n3204), .B(n3110), .Y(n12219) );
  XNOR2X1 U20862 ( .A(n3204), .B(M3_mult_x_15_b_1_), .Y(n12343) );
  XNOR2XL U20863 ( .A(n12265), .B(n11499), .Y(n12220) );
  XNOR2X1 U20864 ( .A(n12282), .B(n3108), .Y(n12232) );
  XNOR2X1 U20865 ( .A(n12282), .B(n3049), .Y(n12223) );
  OAI22XL U20866 ( .A0(n12357), .A1(n12232), .B0(n12284), .B1(n12223), .Y(
        n12239) );
  XNOR2X1 U20867 ( .A(n12265), .B(n12279), .Y(n12236) );
  OAI22XL U20868 ( .A0(n12152), .A1(n12236), .B0(n3185), .B1(n12220), .Y(
        n12238) );
  XNOR2X1 U20869 ( .A(n2980), .B(n3049), .Y(n12245) );
  XNOR2X1 U20870 ( .A(n2980), .B(n3197), .Y(n12227) );
  OAI22XL U20871 ( .A0(n12293), .A1(n12245), .B0(n12227), .B1(n12338), .Y(
        n12244) );
  OAI22XL U20872 ( .A0(n12352), .A1(n11486), .B0(n12222), .B1(n12221), .Y(
        n12243) );
  XNOR2X1 U20873 ( .A(n12282), .B(n3197), .Y(n12356) );
  OAI22XL U20874 ( .A0(n12357), .A1(n12223), .B0(n12284), .B1(n12356), .Y(
        n12366) );
  XNOR2X1 U20875 ( .A(n2980), .B(n5430), .Y(n12226) );
  XNOR2X1 U20876 ( .A(n2980), .B(M3_mult_x_15_b_9_), .Y(n12339) );
  OAI22XL U20877 ( .A0(n12293), .A1(n12226), .B0(n12339), .B1(n12338), .Y(
        n12337) );
  NAND2BXL U20878 ( .AN(n3110), .B(n3204), .Y(n12224) );
  XNOR2X1 U20879 ( .A(n12233), .B(M3_mult_x_15_b_1_), .Y(n12234) );
  OAI22XL U20880 ( .A0(n12352), .A1(n12234), .B0(n12222), .B1(n12228), .Y(
        n12229) );
  OAI22XL U20881 ( .A0(n12357), .A1(n12254), .B0(n12284), .B1(n12232), .Y(
        n12249) );
  XNOR2X1 U20882 ( .A(n12233), .B(n3110), .Y(n12235) );
  OAI22XL U20883 ( .A0(n12352), .A1(n12235), .B0(n12222), .B1(n12234), .Y(
        n12248) );
  XNOR2X1 U20884 ( .A(n12265), .B(n12271), .Y(n12246) );
  CMPR32X1 U20885 ( .A(n12239), .B(n12238), .C(n12237), .CO(n12374), .S(n12240) );
  NOR2XL U20886 ( .A(n12326), .B(n12325), .Y(n12329) );
  CMPR32X1 U20887 ( .A(n12242), .B(n12241), .C(n12240), .CO(n12325), .S(n12324) );
  ADDHXL U20888 ( .A(n12244), .B(n12243), .CO(n12237), .S(n12253) );
  XNOR2X1 U20889 ( .A(n2980), .B(n3108), .Y(n12255) );
  OAI22XL U20890 ( .A0(n12152), .A1(n12266), .B0(n3185), .B1(n12246), .Y(
        n12257) );
  CMPR32X1 U20891 ( .A(n12249), .B(n12248), .C(n12247), .CO(n12241), .S(n12251) );
  NOR2XL U20892 ( .A(n12324), .B(n12323), .Y(n12250) );
  NOR2XL U20893 ( .A(n12329), .B(n12250), .Y(n12332) );
  ADDFHX1 U20894 ( .A(n12253), .B(n12252), .CI(n12251), .CO(n12323), .S(n12317) );
  XNOR2XL U20895 ( .A(n2980), .B(n11499), .Y(n12291) );
  OAI22XL U20896 ( .A0(n12293), .A1(n12291), .B0(n12255), .B1(n12338), .Y(
        n12269) );
  OAI22XL U20897 ( .A0(n12152), .A1(n4002), .B0(n3185), .B1(n12256), .Y(n12268) );
  XNOR2X1 U20898 ( .A(n12265), .B(n3110), .Y(n12267) );
  OAI22XL U20899 ( .A0(n12152), .A1(n12267), .B0(n3185), .B1(n12266), .Y(
        n12304) );
  ADDHXL U20900 ( .A(n12269), .B(n12268), .CO(n12262), .S(n12303) );
  OR2X2 U20901 ( .A(n12315), .B(n12314), .Y(n12270) );
  NAND2XL U20902 ( .A(n12260), .B(n12270), .Y(n12322) );
  XNOR2X1 U20903 ( .A(n2980), .B(n12271), .Y(n12280) );
  INVXL U20904 ( .A(n12275), .Y(n12278) );
  INVXL U20905 ( .A(n12272), .Y(n12273) );
  NAND2XL U20906 ( .A(n11697), .B(n12273), .Y(n12277) );
  NAND2XL U20907 ( .A(n12275), .B(n12274), .Y(n12276) );
  OAI21XL U20908 ( .A0(n12278), .A1(n12277), .B0(n12276), .Y(n12290) );
  XNOR2X1 U20909 ( .A(n2980), .B(n12279), .Y(n12292) );
  AND2XL U20910 ( .A(n12288), .B(n12287), .Y(n12289) );
  AOI21XL U20911 ( .A0(n12290), .A1(n12286), .B0(n12289), .Y(n12302) );
  NOR2BXL U20912 ( .AN(n3110), .B(n3185), .Y(n12308) );
  NOR2XL U20913 ( .A(n12299), .B(n12298), .Y(n12301) );
  NAND2XL U20914 ( .A(n12299), .B(n12298), .Y(n12300) );
  OAI21XL U20915 ( .A0(n12302), .A1(n12301), .B0(n12300), .Y(n12313) );
  CMPR32X1 U20916 ( .A(n12305), .B(n12304), .C(n12303), .CO(n12314), .S(n12311) );
  CMPR32X1 U20917 ( .A(n12308), .B(n12307), .C(n12306), .CO(n12310), .S(n12299) );
  AOI21XL U20918 ( .A0(n12313), .A1(n12309), .B0(n12312), .Y(n12321) );
  AND2X2 U20919 ( .A(n12315), .B(n12314), .Y(n12319) );
  AOI21XL U20920 ( .A0(n12260), .A1(n12319), .B0(n12318), .Y(n12320) );
  OAI21XL U20921 ( .A0(n12322), .A1(n12321), .B0(n12320), .Y(n12331) );
  NAND2XL U20922 ( .A(n12324), .B(n12323), .Y(n12328) );
  NAND2XL U20923 ( .A(n12326), .B(n12325), .Y(n12327) );
  OAI21XL U20924 ( .A0(n12329), .A1(n12328), .B0(n12327), .Y(n12330) );
  AOI21XL U20925 ( .A0(n12332), .A1(n12331), .B0(n12330), .Y(n12384) );
  CMPR32X1 U20926 ( .A(n12335), .B(n12334), .C(n12333), .CO(n12395), .S(n12402) );
  OAI22XL U20927 ( .A0(n12598), .A1(n12343), .B0(n12342), .B1(n12341), .Y(
        n12347) );
  CMPR32X1 U20928 ( .A(n12349), .B(n12348), .C(n12347), .CO(n12393), .S(n12368) );
  OAI22XL U20929 ( .A0(n12352), .A1(n12351), .B0(n12222), .B1(n12350), .Y(
        n12363) );
  OAI22XL U20930 ( .A0(n12357), .A1(n12356), .B0(n12284), .B1(n12355), .Y(
        n12361) );
  CMPR32X1 U20931 ( .A(n12360), .B(n12359), .C(n12358), .CO(n12396), .S(n12391) );
  CMPR32X1 U20932 ( .A(n12375), .B(n12374), .C(n12373), .CO(n12377), .S(n12326) );
  OR2X2 U20933 ( .A(n12378), .B(n12377), .Y(n12376) );
  AND2X2 U20934 ( .A(n12378), .B(n12377), .Y(n12382) );
  AND2X2 U20935 ( .A(n12380), .B(n12379), .Y(n12381) );
  CMPR32X1 U20936 ( .A(n12399), .B(n12398), .C(n12397), .CO(n12405), .S(n12404) );
  NAND2XL U20937 ( .A(n12409), .B(n12408), .Y(n12413) );
  NAND2XL U20938 ( .A(n12411), .B(n12410), .Y(n12412) );
  OAI21XL U20939 ( .A0(n12414), .A1(n12413), .B0(n12412), .Y(n12418) );
  AND2X2 U20940 ( .A(n12416), .B(n12415), .Y(n12417) );
  ADDFHX1 U20941 ( .A(n12435), .B(n12434), .CI(n12433), .CO(n12430), .S(n12465) );
  ADDFHX1 U20942 ( .A(n12441), .B(n12440), .CI(n12439), .CO(n12463), .S(n12471) );
  ADDFHX1 U20943 ( .A(n12450), .B(n12449), .CI(n12448), .CO(n12447), .S(n12459) );
  ADDFHX2 U20944 ( .A(n12471), .B(n12470), .CI(n12469), .CO(n12488), .S(n12428) );
  ADDFHX4 U20945 ( .A(n12479), .B(n12478), .CI(n12477), .CO(n12483), .S(n12485) );
  ADDFHX4 U20946 ( .A(n12487), .B(n12486), .CI(n12485), .CO(n12492), .S(n12491) );
  XNOR2XL U20947 ( .A(n12716), .B(M5_b_18_), .Y(n12527) );
  OAI22XL U20948 ( .A0(n12717), .A1(n12527), .B0(n12718), .B1(n12516), .Y(
        n12533) );
  OAI2BB1XL U20949 ( .A0N(n12523), .A1N(n12597), .B0(M3_a_11_), .Y(n12531) );
  XNOR2X1 U20950 ( .A(n25884), .B(n12803), .Y(n12515) );
  OAI22XL U20951 ( .A0(n12618), .A1(n12534), .B0(n12616), .B1(n12515), .Y(
        n12530) );
  XNOR2X1 U20952 ( .A(n12758), .B(n12701), .Y(n12526) );
  XNOR2X1 U20953 ( .A(n12758), .B(n3198), .Y(n12517) );
  OAI22X1 U20954 ( .A0(n12759), .A1(n12526), .B0(n11749), .B1(n12517), .Y(
        n12529) );
  XNOR2X1 U20955 ( .A(n12732), .B(n3021), .Y(n12524) );
  XNOR2XL U20956 ( .A(n12732), .B(M5_b_18_), .Y(n12546) );
  OAI22XL U20957 ( .A0(n12715), .A1(n12514), .B0(n12746), .B1(n12546), .Y(
        n12545) );
  XNOR2X1 U20958 ( .A(n12758), .B(n3021), .Y(n12540) );
  OAI22XL U20959 ( .A0(n12759), .A1(n12517), .B0(n12760), .B1(n12540), .Y(
        n12538) );
  OAI22XL U20960 ( .A0(n12535), .A1(n12561), .B0(n12995), .B1(n12518), .Y(
        n12520) );
  OAI22XL U20961 ( .A0(n12635), .A1(n12519), .B0(n12633), .B1(
        M3_U3_U1_or2_inv_0__18_), .Y(n12541) );
  CMPR32X1 U20962 ( .A(M4_mult_x_15_n1680), .B(n3190), .C(n12520), .CO(n12537), 
        .S(n12589) );
  OAI22XL U20963 ( .A0(n12597), .A1(n12594), .B0(n12523), .B1(n12522), .Y(
        n12590) );
  OAI22XL U20964 ( .A0(n12715), .A1(n12638), .B0(n12525), .B1(n12524), .Y(
        n12601) );
  XNOR2X1 U20965 ( .A(n12758), .B(n12560), .Y(n12636) );
  OAI22X1 U20966 ( .A0(n12759), .A1(n12636), .B0(n12760), .B1(n12526), .Y(
        n12600) );
  XNOR2X1 U20967 ( .A(n12716), .B(n3201), .Y(n12592) );
  OAI22XL U20968 ( .A0(n12578), .A1(n12592), .B0(n12718), .B1(n12527), .Y(
        n12599) );
  CMPR32X1 U20969 ( .A(n12530), .B(n12529), .C(n12528), .CO(n12585), .S(n12604) );
  CMPR32X1 U20970 ( .A(n12533), .B(n12532), .C(n12531), .CO(n12586), .S(n12603) );
  XNOR2XL U20971 ( .A(n25884), .B(M3_mult_x_15_b_19_), .Y(n12615) );
  OAI22X2 U20972 ( .A0(n12618), .A1(n12615), .B0(n12616), .B1(n12534), .Y(
        n12644) );
  OAI22X1 U20973 ( .A0(n12535), .A1(n16884), .B0(n12995), .B1(n3190), .Y(
        n12619) );
  XNOR2X1 U20974 ( .A(n12716), .B(n12803), .Y(n12555) );
  OAI22XL U20975 ( .A0(n12576), .A1(n12540), .B0(n12760), .B1(n12553), .Y(
        n12557) );
  CMPR32X1 U20976 ( .A(n12545), .B(n12544), .C(n12543), .CO(n12548), .S(n12584) );
  XNOR2XL U20977 ( .A(n12732), .B(M3_mult_x_15_b_19_), .Y(n12554) );
  OAI22XL U20978 ( .A0(n12715), .A1(n12546), .B0(n12746), .B1(n12554), .Y(
        n12564) );
  ADDFHX1 U20979 ( .A(n12549), .B(n12547), .CI(n12548), .CO(n12567), .S(n12550) );
  OAI22XL U20980 ( .A0(n12576), .A1(n12553), .B0(n12760), .B1(n12575), .Y(
        n12573) );
  OAI22XL U20981 ( .A0(n12715), .A1(n12554), .B0(n12746), .B1(n12574), .Y(
        n12572) );
  XNOR2X1 U20982 ( .A(M3_mult_x_15_a_17_), .B(n3202), .Y(n12577) );
  OAI22X1 U20983 ( .A0(n12717), .A1(n12555), .B0(n12718), .B1(n12577), .Y(
        n12571) );
  CMPR32X1 U20984 ( .A(n12561), .B(n12560), .C(n12559), .CO(n12570), .S(n12556) );
  CMPR32X1 U20985 ( .A(n12567), .B(n12566), .C(n12565), .CO(n12777), .S(n12774) );
  CMPR32X1 U20986 ( .A(n12570), .B(n12569), .C(n12568), .CO(n12692), .S(n12581) );
  ADDFHX1 U20987 ( .A(n12573), .B(n12571), .CI(n12572), .CO(n12704), .S(n12583) );
  XNOR2X1 U20988 ( .A(n12732), .B(n12803), .Y(n12699) );
  OAI22XL U20989 ( .A0(n12715), .A1(n12574), .B0(n12746), .B1(n12699), .Y(
        n12698) );
  CMPR32X1 U20990 ( .A(n12586), .B(n12585), .C(n12584), .CO(n12610), .S(n12668) );
  CMPR32X1 U20991 ( .A(n12589), .B(n12588), .C(n12587), .CO(n12606), .S(n12662) );
  CMPR32X1 U20992 ( .A(n18498), .B(n12591), .C(n12590), .CO(n12588), .S(n12627) );
  CMPR32X1 U20993 ( .A(n12604), .B(n12603), .C(n12602), .CO(n12605), .S(n12660) );
  OAI22XL U20994 ( .A0(n12618), .A1(n12617), .B0(n12616), .B1(n12615), .Y(
        n12647) );
  CMPR32X1 U20995 ( .A(n5430), .B(M3_mult_x_15_b_9_), .C(n12619), .CO(n12643), 
        .S(n12646) );
  ADDFHX1 U20996 ( .A(n16965), .B(n12621), .CI(n12620), .CO(n12645), .S(n12623) );
  OAI22XL U20997 ( .A0(n12635), .A1(n12634), .B0(n12633), .B1(n12632), .Y(
        n12642) );
  CMPR32X1 U20998 ( .A(n12647), .B(n12646), .C(n12645), .CO(n12657), .S(n12655) );
  CMPR32X1 U20999 ( .A(n12659), .B(n12658), .C(n12657), .CO(n12671), .S(n12663) );
  ADDFHX1 U21000 ( .A(n12665), .B(n12664), .CI(n12663), .CO(n12669), .S(n12688) );
  ADDFHX4 U21001 ( .A(n12686), .B(n12685), .CI(n12684), .CO(n12766), .S(n12763) );
  INVXL U21002 ( .A(n12985), .Y(n12864) );
  CMPR32X1 U21003 ( .A(n12692), .B(n12691), .C(n12690), .CO(n12782), .S(n12776) );
  CMPR32X1 U21004 ( .A(n12695), .B(n12694), .C(n12693), .CO(n12707), .S(n12702) );
  OAI22XL U21005 ( .A0(n12535), .A1(M3_mult_x_15_b_17_), .B0(n12995), .B1(
        n3196), .Y(n12712) );
  CMPR32X1 U21006 ( .A(n3043), .B(n12712), .C(n12711), .CO(n12734), .S(n12721)
         );
  XNOR2X1 U21007 ( .A(n12758), .B(n12803), .Y(n12729) );
  OAI22XL U21008 ( .A0(n12759), .A1(n12713), .B0(n12760), .B1(n12729), .Y(
        n12728) );
  CMPR32X1 U21009 ( .A(n12728), .B(n12727), .C(n12726), .CO(n12739), .S(n12733) );
  XNOR2X1 U21010 ( .A(n12758), .B(n3202), .Y(n12745) );
  CMPR32X1 U21011 ( .A(n3021), .B(n3201), .C(n12730), .CO(n12743), .S(n12735)
         );
  INVX1 U21012 ( .A(n12736), .Y(n12871) );
  CMPR32X1 U21013 ( .A(n5997), .B(n12741), .C(n12740), .CO(n12749), .S(n12742)
         );
  CMPR32X1 U21014 ( .A(n12744), .B(n12743), .C(n12742), .CO(n12748), .S(n12738) );
  CMPR32X1 U21015 ( .A(n12749), .B(n12748), .C(n12747), .CO(n12792), .S(n12789) );
  CMPR32X1 U21016 ( .A(n3196), .B(M3_mult_x_15_b_19_), .C(n12750), .CO(n12757), 
        .S(n12752) );
  CMPR32X1 U21017 ( .A(n12754), .B(n12753), .C(n12752), .CO(n12755), .S(n12747) );
  CMPR32X1 U21018 ( .A(n12757), .B(n12756), .C(n12755), .CO(n12796), .S(n12791) );
  CMPR32X1 U21019 ( .A(n5960), .B(n12762), .C(n12761), .CO(n12799), .S(n12756)
         );
  NAND2XL U21020 ( .A(n12864), .B(n12984), .Y(n12798) );
  INVXL U21021 ( .A(n12862), .Y(n12771) );
  NAND2XL U21022 ( .A(n12773), .B(n12772), .Y(n12856) );
  NAND2XL U21023 ( .A(n12777), .B(n12776), .Y(n12842) );
  OAI21XL U21024 ( .A0(n12841), .A1(n12849), .B0(n12842), .Y(n12778) );
  NAND2XL U21025 ( .A(n12786), .B(n12785), .Y(n12870) );
  INVXL U21026 ( .A(n12870), .Y(n12787) );
  OAI21XL U21027 ( .A0(n12821), .A1(n12815), .B0(n12822), .Y(n12793) );
  OAI21XL U21028 ( .A0(n12825), .A1(n12829), .B0(n12830), .Y(n12989) );
  CMPR32X1 U21029 ( .A(n12801), .B(n12800), .C(n12799), .CO(n12805), .S(n12795) );
  CMPR32X1 U21030 ( .A(n18673), .B(n12803), .C(n12802), .CO(n12993), .S(n12800) );
  OR2X2 U21031 ( .A(n12805), .B(n12804), .Y(n12988) );
  NAND2X1 U21032 ( .A(n12988), .B(n12986), .Y(n12806) );
  INVXL U21033 ( .A(n12808), .Y(n12809) );
  NAND2XL U21034 ( .A(n12814), .B(n12817), .Y(n12820) );
  INVXL U21035 ( .A(n12824), .Y(n12827) );
  INVXL U21036 ( .A(n12825), .Y(n12826) );
  INVXL U21037 ( .A(n12836), .Y(n12852) );
  AOI21XL U21038 ( .A0(n12852), .A1(n12611), .B0(n12837), .Y(n12838) );
  INVXL U21039 ( .A(n12841), .Y(n12843) );
  NAND2XL U21040 ( .A(n12973), .B(n12977), .Y(n12869) );
  INVXL U21041 ( .A(n12874), .Y(n12876) );
  INVX1 U21042 ( .A(n12930), .Y(n12883) );
  NAND2XL U21043 ( .A(n12925), .B(n12883), .Y(n12885) );
  INVXL U21044 ( .A(n12931), .Y(n12882) );
  INVXL U21045 ( .A(n12886), .Y(n12888) );
  INVXL U21046 ( .A(n12897), .Y(n12899) );
  NAND2XL U21047 ( .A(n12914), .B(n12901), .Y(n12904) );
  INVXL U21048 ( .A(n12902), .Y(n12916) );
  AOI21XL U21049 ( .A0(n12919), .A1(n12901), .B0(n12902), .Y(n12903) );
  NAND2XL U21050 ( .A(n12914), .B(n12893), .Y(n12908) );
  INVXL U21051 ( .A(n12980), .Y(n12912) );
  OAI21XL U21052 ( .A0(n12916), .A1(n12905), .B0(n12915), .Y(n12917) );
  AOI21X1 U21053 ( .A0(n12919), .A1(n12918), .B0(n12917), .Y(n12920) );
  INVXL U21054 ( .A(n12922), .Y(n12924) );
  INVXL U21055 ( .A(n12925), .Y(n12928) );
  INVXL U21056 ( .A(n12926), .Y(n12927) );
  INVXL U21057 ( .A(n12934), .Y(n12935) );
  INVXL U21058 ( .A(n12936), .Y(n12938) );
  NAND2XL U21059 ( .A(n12938), .B(n12937), .Y(n12939) );
  INVX1 U21060 ( .A(M3_U4_U1_enc_tree_2__4__16_), .Y(n18818) );
  INVX1 U21061 ( .A(M3_U4_U1_enc_tree_0__4__16_), .Y(n18840) );
  INVX1 U21062 ( .A(M3_U4_U1_enc_tree_1__4__16_), .Y(n18822) );
  OAI21XL U21063 ( .A0(n12961), .A1(n18818), .B0(n12963), .Y(n12943) );
  OAI21XL U21064 ( .A0(n18797), .A1(M3_U3_U1_enc_tree_2__4__16_), .B0(n12943), 
        .Y(n12948) );
  INVX1 U21065 ( .A(n18800), .Y(n18804) );
  NOR2X1 U21066 ( .A(n13032), .B(n13034), .Y(n12971) );
  INVXL U21067 ( .A(n12981), .Y(n12983) );
  CMPR32X1 U21068 ( .A(n5957), .B(n12994), .C(n12993), .CO(n12998), .S(n12804)
         );
  NOR2X1 U21069 ( .A(n13003), .B(n19024), .Y(n24050) );
  XNOR2X1 U21070 ( .A(n14027), .B(n25860), .Y(n13161) );
  XNOR2X1 U21071 ( .A(n14028), .B(n25860), .Y(n13046) );
  OAI22XL U21072 ( .A0(n13161), .A1(n13721), .B0(n13046), .B1(n13790), .Y(
        n13164) );
  CLKBUFX3 U21073 ( .A(M1_a_1_), .Y(n13769) );
  XNOR2XL U21074 ( .A(n13769), .B(n14030), .Y(n13155) );
  XNOR2XL U21075 ( .A(n13049), .B(n14030), .Y(n13043) );
  AND2X4 U21076 ( .A(n14045), .B(n13041), .Y(n13042) );
  XNOR2X2 U21077 ( .A(M1_b_3_), .B(M1_b_4_), .Y(n13899) );
  XOR2X1 U21078 ( .A(M1_b_4_), .B(n13898), .Y(n13044) );
  XNOR2XL U21079 ( .A(n13769), .B(n4807), .Y(n13064) );
  XOR2X1 U21080 ( .A(M1_b_6_), .B(n4807), .Y(n13048) );
  OAI22XL U21081 ( .A0(n13064), .A1(n13971), .B0(n13053), .B1(n13972), .Y(
        n13067) );
  OAI22XL U21082 ( .A0(n13971), .A1(n13047), .B0(n13050), .B1(n13972), .Y(
        n13073) );
  INVX1 U21083 ( .A(n3214), .Y(n13204) );
  XNOR2XL U21084 ( .A(n14027), .B(n13204), .Y(n13056) );
  AND2X2 U21085 ( .A(n13605), .B(n3181), .Y(n13054) );
  CLKINVX3 U21086 ( .A(n13054), .Y(n13532) );
  XNOR2XL U21087 ( .A(n4565), .B(n13204), .Y(n13055) );
  OAI22X1 U21088 ( .A0(n13157), .A1(n3181), .B0(n13055), .B1(n13532), .Y(
        n13181) );
  XNOR2XL U21089 ( .A(n13863), .B(n4807), .Y(n13160) );
  OAI22XL U21090 ( .A0(n13160), .A1(n13972), .B0(n13053), .B1(n13971), .Y(
        n13158) );
  CLKINVX3 U21091 ( .A(n13054), .Y(n13606) );
  XNOR2X1 U21092 ( .A(n13863), .B(n13844), .Y(n13062) );
  OAI22XL U21093 ( .A0(n13062), .A1(n2997), .B0(n13058), .B1(n13843), .Y(
        n13059) );
  ADDFHX1 U21094 ( .A(n13061), .B(n13060), .CI(n13059), .CO(n13179), .S(n13071) );
  XNOR2XL U21095 ( .A(n13864), .B(n13844), .Y(n13083) );
  OAI22XL U21096 ( .A0(n13062), .A1(n13899), .B0(n13083), .B1(n2997), .Y(
        n13078) );
  XNOR2XL U21097 ( .A(n13049), .B(n4807), .Y(n13063) );
  OAI22XL U21098 ( .A0(n13064), .A1(n13972), .B0(n13063), .B1(n13971), .Y(
        n13077) );
  XNOR2X1 U21099 ( .A(n25865), .B(n25860), .Y(n13074) );
  CMPR32X1 U21100 ( .A(n13068), .B(n13067), .C(n13066), .CO(n13189), .S(n13069) );
  NOR2XL U21101 ( .A(n13148), .B(n13147), .Y(n13151) );
  ADDHXL U21102 ( .A(n13073), .B(n13072), .CO(n13066), .S(n13082) );
  XNOR2X1 U21103 ( .A(n13863), .B(n25860), .Y(n13085) );
  OAI22XL U21104 ( .A0(n13092), .A1(n13606), .B0(n13075), .B1(n3181), .Y(
        n13086) );
  CMPR32X1 U21105 ( .A(n13078), .B(n13077), .C(n13076), .CO(n13070), .S(n13080) );
  NOR2XL U21106 ( .A(n13146), .B(n13145), .Y(n13079) );
  NOR2XL U21107 ( .A(n13151), .B(n13079), .Y(n13154) );
  ADDFHX1 U21108 ( .A(n13082), .B(n13081), .CI(n13080), .CO(n13145), .S(n13138) );
  OAI22XL U21109 ( .A0(n2997), .A1(n13842), .B0(n13084), .B1(n13843), .Y(
        n13096) );
  XNOR2X1 U21110 ( .A(n13864), .B(n25860), .Y(n13115) );
  CMPR32X1 U21111 ( .A(n13088), .B(n13087), .C(n13086), .CO(n13081), .S(n13089) );
  OR2X2 U21112 ( .A(n13138), .B(n13137), .Y(n13141) );
  OAI22XL U21113 ( .A0(n13092), .A1(n3181), .B0(n13113), .B1(n13532), .Y(
        n13126) );
  ADDHXL U21114 ( .A(n13096), .B(n13095), .CO(n13090), .S(n13124) );
  OR2X2 U21115 ( .A(n13136), .B(n13135), .Y(n13097) );
  NAND2XL U21116 ( .A(n13141), .B(n13097), .Y(n13144) );
  XNOR2XL U21117 ( .A(n13864), .B(n13204), .Y(n13107) );
  OAI22XL U21118 ( .A0(n13769), .A1(n13606), .B0(n13107), .B1(n3181), .Y(
        n13102) );
  INVXL U21119 ( .A(n13102), .Y(n13105) );
  INVXL U21120 ( .A(n13098), .Y(n13099) );
  NAND2XL U21121 ( .A(n13100), .B(n13099), .Y(n13104) );
  NAND2XL U21122 ( .A(n13102), .B(n13101), .Y(n13103) );
  OAI21XL U21123 ( .A0(n13105), .A1(n13104), .B0(n13103), .Y(n13112) );
  XNOR2XL U21124 ( .A(n13863), .B(n13204), .Y(n13114) );
  AOI21XL U21125 ( .A0(n13112), .A1(n13109), .B0(n6204), .Y(n13123) );
  OAI22XL U21126 ( .A0(n13114), .A1(n13606), .B0(n13113), .B1(n3181), .Y(
        n13128) );
  NOR2XL U21127 ( .A(n13120), .B(n13119), .Y(n13122) );
  NAND2XL U21128 ( .A(n13120), .B(n13119), .Y(n13121) );
  OAI21XL U21129 ( .A0(n13123), .A1(n13122), .B0(n13121), .Y(n13134) );
  CMPR32X1 U21130 ( .A(n13126), .B(n13125), .C(n13124), .CO(n13135), .S(n13131) );
  CMPR32X1 U21131 ( .A(n13129), .B(n13128), .C(n13127), .CO(n13130), .S(n13120) );
  OR2XL U21132 ( .A(n13131), .B(n13130), .Y(n13133) );
  AOI21XL U21133 ( .A0(n13134), .A1(n13133), .B0(n13132), .Y(n13143) );
  AND2X2 U21134 ( .A(n13138), .B(n13137), .Y(n13139) );
  AOI21XL U21135 ( .A0(n13141), .A1(n13140), .B0(n13139), .Y(n13142) );
  OAI21XL U21136 ( .A0(n13144), .A1(n13143), .B0(n13142), .Y(n13153) );
  NAND2XL U21137 ( .A(n13146), .B(n13145), .Y(n13150) );
  NAND2XL U21138 ( .A(n13148), .B(n13147), .Y(n13149) );
  OAI21XL U21139 ( .A0(n13151), .A1(n13150), .B0(n13149), .Y(n13152) );
  AOI21XL U21140 ( .A0(n13154), .A1(n13153), .B0(n13152), .Y(n13201) );
  XNOR2XL U21141 ( .A(n13864), .B(n14030), .Y(n13171) );
  OAI22XL U21142 ( .A0(n13156), .A1(n2997), .B0(n13168), .B1(n13843), .Y(
        n13177) );
  XNOR2XL U21143 ( .A(n14118), .B(n13204), .Y(n13175) );
  OAI22XL U21144 ( .A0(n13157), .A1(n13606), .B0(n13175), .B1(n3181), .Y(
        n13176) );
  ADDHXL U21145 ( .A(n13159), .B(n13158), .CO(n13184), .S(n13180) );
  NOR2BX1 U21146 ( .AN(n13049), .B(n3173), .Y(n13167) );
  XNOR2XL U21147 ( .A(n25865), .B(n4807), .Y(n13172) );
  XNOR2X1 U21148 ( .A(n4565), .B(n25860), .Y(n13170) );
  OAI22XL U21149 ( .A0(n13161), .A1(n13790), .B0(n13170), .B1(n13721), .Y(
        n13165) );
  ADDFHX1 U21150 ( .A(n13164), .B(n13163), .CI(n13162), .CO(n13182), .S(n13190) );
  ADDFHX1 U21151 ( .A(n13167), .B(n13166), .CI(n13165), .CO(n13236), .S(n13183) );
  OAI22X1 U21152 ( .A0(n13206), .A1(n13899), .B0(n13168), .B1(n2997), .Y(
        n13211) );
  XNOR2XL U21153 ( .A(n13769), .B(M1_b_11_), .Y(n13225) );
  XNOR2XL U21154 ( .A(M1_a_0_), .B(M1_b_11_), .Y(n13169) );
  XNOR2XL U21155 ( .A(n13863), .B(n14030), .Y(n13207) );
  XNOR2XL U21156 ( .A(n13919), .B(n4807), .Y(n13209) );
  NAND2BXL U21157 ( .AN(n13049), .B(n25861), .Y(n13174) );
  OAI22XL U21158 ( .A0(n14080), .A1(n5489), .B0(n13174), .B1(n3173), .Y(n13227) );
  BUFX3 U21159 ( .A(M1_a_11_), .Y(n14117) );
  XNOR2XL U21160 ( .A(n14117), .B(n13204), .Y(n13205) );
  OAI22XL U21161 ( .A0(n13205), .A1(n3181), .B0(n13175), .B1(n13532), .Y(
        n13226) );
  CMPR32X1 U21162 ( .A(n13178), .B(n13177), .C(n13176), .CO(n13245), .S(n13187) );
  ADDFHX1 U21163 ( .A(n13180), .B(n13181), .CI(n13179), .CO(n13186), .S(n13188) );
  ADDFHX1 U21164 ( .A(n13184), .B(n13183), .CI(n13182), .CO(n13244), .S(n13185) );
  OR2X2 U21165 ( .A(n13195), .B(n13194), .Y(n13198) );
  ADDFHX1 U21166 ( .A(n13187), .B(n13186), .CI(n13185), .CO(n13194), .S(n13193) );
  CMPR32X1 U21167 ( .A(n13190), .B(n13189), .C(n13188), .CO(n13192), .S(n13148) );
  OR2X2 U21168 ( .A(n13193), .B(n13192), .Y(n13191) );
  AND2XL U21169 ( .A(n13193), .B(n13192), .Y(n13197) );
  AOI21XL U21170 ( .A0(n13198), .A1(n13197), .B0(n13196), .Y(n13199) );
  OAI21XL U21171 ( .A0(n13201), .A1(n13200), .B0(n13199), .Y(n13256) );
  OAI22XL U21172 ( .A0(n14121), .A1(n14119), .B0(n13202), .B1(n14120), .Y(
        n13264) );
  XNOR2XL U21173 ( .A(n13863), .B(n25861), .Y(n13284) );
  XNOR2XL U21174 ( .A(n13864), .B(n25861), .Y(n13224) );
  XNOR2XL U21175 ( .A(n14196), .B(n13204), .Y(n13222) );
  OAI22XL U21176 ( .A0(n13205), .A1(n13606), .B0(n13222), .B1(n3181), .Y(
        n13229) );
  OAI22XL U21177 ( .A0(n13206), .A1(n2997), .B0(n13220), .B1(n13843), .Y(
        n13228) );
  XNOR2XL U21178 ( .A(n25865), .B(n14030), .Y(n13219) );
  OAI22XL U21179 ( .A0(n13207), .A1(n14044), .B0(n13219), .B1(n13974), .Y(
        n13217) );
  XNOR2X1 U21180 ( .A(n14118), .B(n13693), .Y(n13218) );
  XNOR2XL U21181 ( .A(n14028), .B(n4807), .Y(n13221) );
  OAI22XL U21182 ( .A0(n13209), .A1(n13971), .B0(n13221), .B1(n13972), .Y(
        n13215) );
  XNOR2XL U21183 ( .A(n13919), .B(n14030), .Y(n13266) );
  XNOR2XL U21184 ( .A(n14027), .B(n4807), .Y(n13257) );
  BUFX3 U21185 ( .A(M1_a_13_), .Y(n14195) );
  XNOR2XL U21186 ( .A(n14195), .B(n13605), .Y(n13260) );
  OAI22XL U21187 ( .A0(n13260), .A1(n3181), .B0(n13222), .B1(n13532), .Y(
        n13269) );
  XNOR2XL U21188 ( .A(n13049), .B(n14156), .Y(n13223) );
  OAI22XL U21189 ( .A0(n13259), .A1(n14120), .B0(n13223), .B1(n14121), .Y(
        n13268) );
  OAI22X1 U21190 ( .A0(n13225), .A1(n14080), .B0(n13224), .B1(n3173), .Y(
        n13233) );
  ADDHXL U21191 ( .A(n13227), .B(n13226), .CO(n13232), .S(n13212) );
  CMPR32X1 U21192 ( .A(n13230), .B(n13229), .C(n13228), .CO(n13275), .S(n13231) );
  NOR2X1 U21193 ( .A(n13250), .B(n13249), .Y(n13253) );
  CMPR32X1 U21194 ( .A(n13242), .B(n13241), .C(n13240), .CO(n13249), .S(n13248) );
  CMPR32X1 U21195 ( .A(n13245), .B(n13244), .C(n13243), .CO(n13247), .S(n13195) );
  NOR2XL U21196 ( .A(n13248), .B(n13247), .Y(n13246) );
  NOR2XL U21197 ( .A(n13253), .B(n13246), .Y(n13255) );
  NAND2XL U21198 ( .A(n13248), .B(n13247), .Y(n13252) );
  NAND2XL U21199 ( .A(n13250), .B(n13249), .Y(n13251) );
  OAI21XL U21200 ( .A0(n13253), .A1(n13252), .B0(n13251), .Y(n13254) );
  AOI21XL U21201 ( .A0(n13256), .A1(n13255), .B0(n13254), .Y(n13354) );
  XNOR2XL U21202 ( .A(n4565), .B(n4807), .Y(n13278) );
  OAI22XL U21203 ( .A0(n13257), .A1(n13971), .B0(n13278), .B1(n13972), .Y(
        n13295) );
  XNOR2XL U21204 ( .A(n13864), .B(n14156), .Y(n13279) );
  OAI22XL U21205 ( .A0(n13260), .A1(n13606), .B0(n13282), .B1(n3181), .Y(
        n13293) );
  XNOR2XL U21206 ( .A(n14027), .B(n14030), .Y(n13329) );
  XNOR2XL U21207 ( .A(n14028), .B(n14030), .Y(n13265) );
  OAI22XL U21208 ( .A0(n13329), .A1(n14029), .B0(n13265), .B1(n14044), .Y(
        n13332) );
  XOR2X1 U21209 ( .A(M1_b_14_), .B(n25862), .Y(n13261) );
  OAI22X1 U21210 ( .A0(n13316), .A1(n14198), .B0(n13262), .B1(n14208), .Y(
        n13331) );
  XNOR2X1 U21211 ( .A(n14196), .B(n25860), .Y(n13285) );
  ADDHXL U21212 ( .A(n13264), .B(n13263), .CO(n13273), .S(n13276) );
  OAI22XL U21213 ( .A0(n13266), .A1(n14044), .B0(n13265), .B1(n13974), .Y(
        n13272) );
  OAI22XL U21214 ( .A0(n13267), .A1(n2997), .B0(n13277), .B1(n13843), .Y(
        n13271) );
  CMPR32X1 U21215 ( .A(n13270), .B(n13269), .C(n13268), .CO(n13304), .S(n13300) );
  CMPR32X1 U21216 ( .A(n13271), .B(n13272), .C(n13273), .CO(n13333), .S(n13303) );
  ADDFHX1 U21217 ( .A(n13276), .B(n13275), .CI(n13274), .CO(n13302), .S(n13310) );
  OAI22XL U21218 ( .A0(n13314), .A1(n13899), .B0(n13277), .B1(n2997), .Y(
        n13313) );
  XNOR2XL U21219 ( .A(n4567), .B(n4807), .Y(n13319) );
  OAI22X1 U21220 ( .A0(n13319), .A1(n13972), .B0(n13278), .B1(n13971), .Y(
        n13312) );
  BUFX3 U21221 ( .A(M1_a_15_), .Y(n14235) );
  XNOR2XL U21222 ( .A(n14235), .B(n13605), .Y(n13328) );
  NOR2BX1 U21223 ( .AN(n13049), .B(n14198), .Y(n13289) );
  OAI22XL U21224 ( .A0(n13286), .A1(n13790), .B0(n13285), .B1(n13721), .Y(
        n13287) );
  ADDFHX1 U21225 ( .A(n13289), .B(n13288), .CI(n13287), .CO(n13323), .S(n13298) );
  ADDFHX1 U21226 ( .A(n13292), .B(n13291), .CI(n13290), .CO(n13297), .S(n13301) );
  ADDFHX1 U21227 ( .A(n13295), .B(n13294), .CI(n13293), .CO(n13335), .S(n13296) );
  ADDFHX1 U21228 ( .A(n13298), .B(n13297), .CI(n13296), .CO(n13320), .S(n13307) );
  ADDFHX1 U21229 ( .A(n13313), .B(n13312), .CI(n13311), .CO(n13383), .S(n13322) );
  XNOR2XL U21230 ( .A(n14196), .B(n4848), .Y(n13392) );
  OAI22XL U21231 ( .A0(n13314), .A1(n2997), .B0(n13392), .B1(n13843), .Y(
        n13377) );
  XNOR2XL U21232 ( .A(n14236), .B(M1_b_3_), .Y(n13390) );
  OAI22XL U21233 ( .A0(n13317), .A1(n14157), .B0(n13359), .B1(n14120), .Y(
        n13389) );
  XNOR2XL U21234 ( .A(n14028), .B(M1_b_11_), .Y(n13360) );
  OAI22X1 U21235 ( .A0(n13318), .A1(n14080), .B0(n13360), .B1(n3173), .Y(
        n13388) );
  XNOR2XL U21236 ( .A(n14118), .B(n4807), .Y(n13355) );
  OAI22XL U21237 ( .A0(n13319), .A1(n13971), .B0(n13355), .B1(n13972), .Y(
        n13387) );
  ADDFHX1 U21238 ( .A(n13325), .B(n13324), .CI(n13323), .CO(n13410), .S(n13321) );
  CMPR22X1 U21239 ( .A(n13327), .B(n13326), .CO(n13371), .S(n13324) );
  XNOR2XL U21240 ( .A(n4565), .B(n14030), .Y(n13361) );
  OAI22XL U21241 ( .A0(n13329), .A1(n14044), .B0(n13361), .B1(n13974), .Y(
        n13372) );
  ADDFHX1 U21242 ( .A(n13332), .B(n13331), .CI(n13330), .CO(n13369), .S(n13334) );
  ADDFHX1 U21243 ( .A(n13335), .B(n13334), .CI(n13333), .CO(n13408), .S(n13338) );
  NAND2XL U21244 ( .A(n13339), .B(n13350), .Y(n13353) );
  NAND2XL U21245 ( .A(n13341), .B(n13340), .Y(n13345) );
  NAND2XL U21246 ( .A(n13343), .B(n13342), .Y(n13344) );
  AND2X2 U21247 ( .A(n13348), .B(n13347), .Y(n13349) );
  OAI21XL U21248 ( .A0(n13354), .A1(n13353), .B0(n13352), .Y(n13469) );
  XNOR2XL U21249 ( .A(n14117), .B(n4807), .Y(n13368) );
  OAI22XL U21250 ( .A0(n13368), .A1(n13972), .B0(n13355), .B1(n13971), .Y(
        n13395) );
  XNOR2XL U21251 ( .A(n13049), .B(n14228), .Y(n13358) );
  NAND2X4 U21252 ( .A(n13357), .B(n14250), .Y(n14249) );
  OAI22XL U21253 ( .A0(n13403), .A1(n14227), .B0(n13358), .B1(n14249), .Y(
        n13394) );
  XNOR2XL U21254 ( .A(n13919), .B(n14156), .Y(n13401) );
  XNOR2XL U21255 ( .A(n14027), .B(M1_b_11_), .Y(n13402) );
  OAI22XL U21256 ( .A0(n13402), .A1(n3173), .B0(n13360), .B1(n14080), .Y(
        n13380) );
  XNOR2XL U21257 ( .A(n4567), .B(n14030), .Y(n13364) );
  OAI22X1 U21258 ( .A0(n13364), .A1(n14029), .B0(n13361), .B1(n14044), .Y(
        n13379) );
  CLKINVX3 U21259 ( .A(n13428), .Y(n14268) );
  XNOR2XL U21260 ( .A(n25865), .B(n25862), .Y(n13448) );
  XNOR2XL U21261 ( .A(n14196), .B(n4807), .Y(n13451) );
  OAI22XL U21262 ( .A0(n13368), .A1(n13971), .B0(n13451), .B1(n13972), .Y(
        n13431) );
  CMPR32X1 U21263 ( .A(n13380), .B(n13379), .C(n13378), .CO(n13453), .S(n13384) );
  ADDFHX1 U21264 ( .A(n13383), .B(n13382), .CI(n13381), .CO(n13411), .S(n13419) );
  ADDFHX1 U21265 ( .A(n13389), .B(n13388), .CI(n13387), .CO(n13407), .S(n13381) );
  BUFX3 U21266 ( .A(M1_a_17_), .Y(n14265) );
  XNOR2XL U21267 ( .A(n14265), .B(n13605), .Y(n13404) );
  OAI22XL U21268 ( .A0(n13404), .A1(n3181), .B0(n13391), .B1(n13532), .Y(
        n13397) );
  XNOR2X1 U21269 ( .A(n14195), .B(n4848), .Y(n13400) );
  OAI22XL U21270 ( .A0(n13400), .A1(n13899), .B0(n13392), .B1(n2997), .Y(
        n13396) );
  OAI22X1 U21271 ( .A0(n13400), .A1(n2997), .B0(n13446), .B1(n13843), .Y(
        n13444) );
  OAI22XL U21272 ( .A0(n13401), .A1(n14157), .B0(n13449), .B1(n14120), .Y(
        n13443) );
  XNOR2XL U21273 ( .A(n4565), .B(n25861), .Y(n13423) );
  OAI22XL U21274 ( .A0(n13402), .A1(n14080), .B0(n13423), .B1(n3173), .Y(
        n13436) );
  XNOR2XL U21275 ( .A(n13864), .B(n14228), .Y(n13422) );
  OAI22XL U21276 ( .A0(n13404), .A1(n13606), .B0(n13430), .B1(n3181), .Y(
        n13434) );
  ADDFHX4 U21277 ( .A(n13407), .B(n13406), .CI(n13405), .CO(n13438), .S(n13416) );
  ADDFHX1 U21278 ( .A(n13410), .B(n13409), .CI(n13408), .CO(n13415), .S(n13417) );
  ADDFHX4 U21279 ( .A(n13413), .B(n13412), .CI(n13411), .CO(n13456), .S(n13414) );
  ADDFHX1 U21280 ( .A(n13416), .B(n13415), .CI(n13414), .CO(n13461), .S(n13460) );
  OR2X2 U21281 ( .A(n13460), .B(n13459), .Y(n13420) );
  NAND2XL U21282 ( .A(n13420), .B(n13463), .Y(n13458) );
  XNOR2XL U21283 ( .A(n13863), .B(n14228), .Y(n13496) );
  XNOR2XL U21284 ( .A(n4567), .B(n25861), .Y(n13497) );
  OAI22XL U21285 ( .A0(n13497), .A1(n3173), .B0(n13423), .B1(n14080), .Y(
        n13478) );
  XNOR2XL U21286 ( .A(n14288), .B(n13605), .Y(n13476) );
  ADDFHX1 U21287 ( .A(n13433), .B(n13432), .CI(n13431), .CO(n13474), .S(n13424) );
  XNOR2XL U21288 ( .A(n13769), .B(n25863), .Y(n13494) );
  XNOR2XL U21289 ( .A(n13049), .B(n25863), .Y(n13447) );
  OAI22X1 U21290 ( .A0(n13494), .A1(n14268), .B0(n13447), .B1(n14282), .Y(
        n13491) );
  OAI22XL U21291 ( .A0(n13483), .A1(n14198), .B0(n13448), .B1(n14208), .Y(
        n13490) );
  XNOR2XL U21292 ( .A(n14027), .B(n14156), .Y(n13495) );
  OAI22XL U21293 ( .A0(n13495), .A1(n14120), .B0(n13449), .B1(n14121), .Y(
        n13472) );
  XNOR2XL U21294 ( .A(n14195), .B(n4807), .Y(n13493) );
  NOR2XL U21295 ( .A(n13465), .B(n13464), .Y(n13466) );
  NOR2XL U21296 ( .A(n13458), .B(n13466), .Y(n13468) );
  ADDFHX1 U21297 ( .A(n13475), .B(n13474), .CI(n13473), .CO(n13545), .S(n13500) );
  XNOR2X2 U21298 ( .A(M1_b_20_), .B(M1_b_19_), .Y(n14291) );
  OAI22X1 U21299 ( .A0(n13476), .A1(n13606), .B0(n13533), .B1(n3181), .Y(
        n13514) );
  XNOR2XL U21300 ( .A(n14266), .B(n4848), .Y(n13534) );
  OAI22XL U21301 ( .A0(n13477), .A1(n2997), .B0(n13534), .B1(n13843), .Y(
        n13513) );
  OAI22XL U21302 ( .A0(n13481), .A1(n14044), .B0(n13540), .B1(n13974), .Y(
        n13527) );
  XNOR2XL U21303 ( .A(n25864), .B(n13693), .Y(n13538) );
  OAI22XL U21304 ( .A0(n13483), .A1(n14208), .B0(n13541), .B1(n14198), .Y(
        n13525) );
  ADDFHX1 U21305 ( .A(n13492), .B(n13491), .CI(n13490), .CO(n13521), .S(n13488) );
  XNOR2XL U21306 ( .A(n14236), .B(n4807), .Y(n13506) );
  XNOR2XL U21307 ( .A(n13864), .B(n25863), .Y(n13512) );
  OAI22X1 U21308 ( .A0(n13494), .A1(n14282), .B0(n13512), .B1(n14251), .Y(
        n13536) );
  XNOR2XL U21309 ( .A(M1_a_8_), .B(n14156), .Y(n13539) );
  OAI22XL U21310 ( .A0(n13495), .A1(n14157), .B0(n13539), .B1(n14120), .Y(
        n13535) );
  XNOR2XL U21311 ( .A(n25865), .B(n14228), .Y(n13543) );
  OAI22XL U21312 ( .A0(n13496), .A1(n14249), .B0(n13543), .B1(n14250), .Y(
        n13530) );
  XNOR2XL U21313 ( .A(n14118), .B(n25861), .Y(n13531) );
  OAI22XL U21314 ( .A0(n13497), .A1(n14080), .B0(n13531), .B1(n3173), .Y(
        n13529) );
  ADDFHX1 U21315 ( .A(n13505), .B(n13504), .CI(n13503), .CO(n13590), .S(n13465) );
  XNOR2XL U21316 ( .A(n14235), .B(n4807), .Y(n13563) );
  OAI22XL U21317 ( .A0(n13563), .A1(n13972), .B0(n13506), .B1(n13971), .Y(
        n13580) );
  NAND2X2 U21318 ( .A(n3229), .B(w1[149]), .Y(n13508) );
  XOR2X1 U21319 ( .A(n23173), .B(M1_b_20_), .Y(n13509) );
  XNOR2XL U21320 ( .A(n13863), .B(n25863), .Y(n13555) );
  ADDFHX1 U21321 ( .A(n13515), .B(n13514), .CI(n13513), .CO(n13578), .S(n13518) );
  XNOR2XL U21322 ( .A(n14117), .B(M1_b_11_), .Y(n13575) );
  OAI22XL U21323 ( .A0(n13575), .A1(n3173), .B0(n13531), .B1(n14080), .Y(
        n13554) );
  BUFX3 U21324 ( .A(M1_a_21_), .Y(n14306) );
  XNOR2XL U21325 ( .A(n14306), .B(n13605), .Y(n13564) );
  OAI22XL U21326 ( .A0(n13565), .A1(n13899), .B0(n13534), .B1(n2997), .Y(
        n13552) );
  ADDFHX1 U21327 ( .A(n13537), .B(n13536), .CI(n13535), .CO(n13559), .S(n13520) );
  XNOR2XL U21328 ( .A(n4567), .B(n14156), .Y(n13576) );
  XNOR2XL U21329 ( .A(n14195), .B(n14030), .Y(n13577) );
  OAI22XL U21330 ( .A0(n13577), .A1(n14029), .B0(n13540), .B1(n14044), .Y(
        n13572) );
  OAI22XL U21331 ( .A0(n13566), .A1(n14198), .B0(n13541), .B1(n14208), .Y(
        n13562) );
  XNOR2XL U21332 ( .A(n13769), .B(n23173), .Y(n13567) );
  XNOR2XL U21333 ( .A(M1_a_0_), .B(n23173), .Y(n13542) );
  XNOR2XL U21334 ( .A(n13919), .B(n14228), .Y(n13568) );
  OAI22XL U21335 ( .A0(n13568), .A1(n14227), .B0(n13543), .B1(n14249), .Y(
        n13560) );
  XNOR2X1 U21336 ( .A(M1_a_4_), .B(n25863), .Y(n13621) );
  XNOR2X1 U21337 ( .A(n14307), .B(n13693), .Y(n13620) );
  OAI22XL U21338 ( .A0(n13556), .A1(n13790), .B0(n13620), .B1(n13721), .Y(
        n13597) );
  XOR3X2 U21339 ( .A(n13635), .B(n13634), .C(n13636), .Y(n13627) );
  XNOR2XL U21340 ( .A(n14266), .B(n4807), .Y(n13617) );
  OAI22XL U21341 ( .A0(n13563), .A1(n13971), .B0(n13617), .B1(n13972), .Y(
        n13615) );
  OAI22XL U21342 ( .A0(n13564), .A1(n13606), .B0(n13607), .B1(n3181), .Y(
        n13614) );
  OAI22XL U21343 ( .A0(n13565), .A1(n2997), .B0(n13601), .B1(n13843), .Y(
        n13613) );
  XNOR2XL U21344 ( .A(M1_a_8_), .B(M1_b_15_), .Y(n13618) );
  OAI22XL U21345 ( .A0(n13566), .A1(n14208), .B0(n13618), .B1(n14198), .Y(
        n13630) );
  XNOR2XL U21346 ( .A(n13864), .B(n23173), .Y(n13603) );
  ADDFHX1 U21347 ( .A(n13571), .B(n13570), .CI(n13569), .CO(n13624), .S(n13586) );
  XNOR2XL U21348 ( .A(n14196), .B(M1_b_11_), .Y(n13608) );
  OAI22XL U21349 ( .A0(n13575), .A1(n14080), .B0(n13608), .B1(n3173), .Y(
        n13633) );
  XNOR2XL U21350 ( .A(n14118), .B(n14156), .Y(n13619) );
  OAI22XL U21351 ( .A0(n13577), .A1(n14044), .B0(n13600), .B1(n13974), .Y(
        n13631) );
  ADDFHX1 U21352 ( .A(n13580), .B(n13579), .CI(n13578), .CO(n13639), .S(n13583) );
  ADDFHX1 U21353 ( .A(n13583), .B(n13582), .CI(n13581), .CO(n13622), .S(n13589) );
  CMPR32X1 U21354 ( .A(n13586), .B(n13585), .C(n13584), .CO(n13642), .S(n13587) );
  ADDFHX1 U21355 ( .A(n13599), .B(n13598), .CI(n13597), .CO(n13686), .S(n13636) );
  XNOR2X1 U21356 ( .A(n14288), .B(n4848), .Y(n13652) );
  OAI22X1 U21357 ( .A0(n13652), .A1(n13899), .B0(n13601), .B1(n2997), .Y(
        n13665) );
  XNOR2XL U21358 ( .A(n13863), .B(n23173), .Y(n13677) );
  OAI22XL U21359 ( .A0(n13607), .A1(n13606), .B0(n3181), .B1(n13605), .Y(
        n13657) );
  XNOR2XL U21360 ( .A(n14195), .B(n25861), .Y(n13667) );
  OAI22XL U21361 ( .A0(n13667), .A1(n3173), .B0(n13608), .B1(n14080), .Y(
        n13656) );
  CLKINVX3 U21362 ( .A(n14353), .Y(n14289) );
  OAI21XL U21363 ( .A0(n14289), .A1(n13049), .B0(n2993), .Y(n13669) );
  OAI22XL U21364 ( .A0(n2993), .A1(n13049), .B0(n14356), .B1(n13769), .Y(
        n13668) );
  CMPR32X1 U21365 ( .A(n13615), .B(n13614), .C(n13613), .CO(n13747), .S(n13611) );
  XNOR2XL U21366 ( .A(n14027), .B(n14228), .Y(n13649) );
  XNOR2XL U21367 ( .A(n14265), .B(n4807), .Y(n13654) );
  XNOR2XL U21368 ( .A(n14117), .B(n14156), .Y(n13666) );
  XNOR2XL U21369 ( .A(n13919), .B(M1_b_19_), .Y(n13651) );
  OAI22XL U21370 ( .A0(n13651), .A1(n14268), .B0(n13621), .B1(n14282), .Y(
        n13658) );
  ADDFHX2 U21371 ( .A(n13624), .B(n13623), .CI(n13622), .CO(n13816), .S(n13643) );
  OAI21XL U21372 ( .A0(n13636), .A1(n13635), .B0(n13634), .Y(n13638) );
  NAND2XL U21373 ( .A(n13636), .B(n13635), .Y(n13637) );
  NAND2X1 U21374 ( .A(n13638), .B(n13637), .Y(n13708) );
  ADDFHX2 U21375 ( .A(n13644), .B(n13643), .CI(n13642), .CO(n13645), .S(n13596) );
  OAI22XL U21376 ( .A0(n13651), .A1(n14282), .B0(n13690), .B1(n14251), .Y(
        n13687) );
  XNOR2X1 U21377 ( .A(n14307), .B(n4848), .Y(n13701) );
  XNOR2XL U21378 ( .A(n25864), .B(n4807), .Y(n13697) );
  OAI22XL U21379 ( .A0(n13654), .A1(n13971), .B0(n13697), .B1(n13972), .Y(
        n13673) );
  CMPR32X1 U21380 ( .A(n13657), .B(n13656), .C(n13655), .CO(n13702), .S(n13684) );
  OR2X2 U21381 ( .A(n13664), .B(n13665), .Y(n13662) );
  OAI22XL U21382 ( .A0(n13666), .A1(n14157), .B0(n13698), .B1(n14120), .Y(
        n13672) );
  OAI22XL U21383 ( .A0(n13667), .A1(n14080), .B0(n13695), .B1(n3173), .Y(
        n13671) );
  ADDHXL U21384 ( .A(n13669), .B(n13668), .CO(n13670), .S(n13655) );
  ADDFHX1 U21385 ( .A(n13672), .B(n4762), .CI(n13670), .CO(n13741), .S(n13705)
         );
  XNOR2XL U21386 ( .A(n25865), .B(n23173), .Y(n13696) );
  OAI22XL U21387 ( .A0(n13677), .A1(n6191), .B0(n13696), .B1(n14298), .Y(
        n13682) );
  OAI22X1 U21388 ( .A0(n2993), .A1(n13769), .B0(n14356), .B1(n13864), .Y(
        n13692) );
  ADDFHX1 U21389 ( .A(n13689), .B(n13688), .CI(n13687), .CO(n13713), .S(n13704) );
  OAI22XL U21390 ( .A0(n13737), .A1(n14268), .B0(n13690), .B1(n14282), .Y(
        n13719) );
  CMPR32X1 U21391 ( .A(n13049), .B(n13692), .C(n13691), .CO(n13718), .S(n13681) );
  XNOR2XL U21392 ( .A(n13919), .B(n23173), .Y(n13723) );
  XNOR2XL U21393 ( .A(n14288), .B(n4807), .Y(n13727) );
  OAI22XL U21394 ( .A0(n13727), .A1(n13972), .B0(n13697), .B1(n13971), .Y(
        n13726) );
  XNOR2XL U21395 ( .A(n14195), .B(n14156), .Y(n13728) );
  XNOR2XL U21396 ( .A(n14265), .B(n14030), .Y(n13729) );
  OAI22XL U21397 ( .A0(n13729), .A1(n14029), .B0(n13699), .B1(n14044), .Y(
        n13724) );
  XNOR2XL U21398 ( .A(n14117), .B(M1_b_15_), .Y(n13722) );
  OAI22X1 U21399 ( .A0(n13722), .A1(n14198), .B0(n13700), .B1(n14208), .Y(
        n13735) );
  XNOR2X1 U21400 ( .A(n14306), .B(n4848), .Y(n13736) );
  OAI22X2 U21401 ( .A0(n13736), .A1(n13899), .B0(n13701), .B1(n2997), .Y(
        n13734) );
  XNOR2XL U21402 ( .A(n4567), .B(n14228), .Y(n13738) );
  CMPR32X1 U21403 ( .A(n13710), .B(n13709), .C(n13708), .CO(n13803), .S(n13810) );
  OAI22XL U21404 ( .A0(n2993), .A1(n13863), .B0(n14356), .B1(n25865), .Y(
        n13767) );
  CMPR32X1 U21405 ( .A(n13100), .B(n13716), .C(n13715), .CO(n13770), .S(n13717) );
  XNOR2XL U21406 ( .A(n14196), .B(M1_b_15_), .Y(n13781) );
  OAI22X1 U21407 ( .A0(n13722), .A1(n14208), .B0(n13781), .B1(n14198), .Y(
        n13774) );
  XNOR2XL U21408 ( .A(n14028), .B(n23173), .Y(n13780) );
  OAI22XL U21409 ( .A0(n13723), .A1(n6191), .B0(n13780), .B1(n14298), .Y(
        n13773) );
  XNOR2XL U21410 ( .A(n14307), .B(n4807), .Y(n13777) );
  XNOR2XL U21411 ( .A(n14236), .B(n14156), .Y(n13792) );
  XNOR2XL U21412 ( .A(n25864), .B(n14030), .Y(n13779) );
  OAI22XL U21413 ( .A0(n13736), .A1(n2997), .B0(n13776), .B1(n13843), .Y(
        n13799) );
  XNOR2XL U21414 ( .A(n4565), .B(n25863), .Y(n13778) );
  XNOR2X1 U21415 ( .A(n14118), .B(n14228), .Y(n13766) );
  OAI22XL U21416 ( .A0(n13738), .A1(n14249), .B0(n13766), .B1(n14250), .Y(
        n13797) );
  XOR3X2 U21417 ( .A(n13786), .B(n13787), .C(n13785), .Y(n13758) );
  ADDFHX1 U21418 ( .A(n13741), .B(n13740), .CI(n13739), .CO(n13757), .S(n13742) );
  ADDFHX1 U21419 ( .A(n13747), .B(n13746), .CI(n13745), .CO(n13814), .S(n13751) );
  ADDFHX4 U21420 ( .A(n13762), .B(n13761), .CI(n13760), .CO(n13825), .S(n13800) );
  XNOR2XL U21421 ( .A(n14117), .B(n14228), .Y(n13839) );
  CMPR32X1 U21422 ( .A(n13769), .B(n13768), .C(n13767), .CO(n13866), .S(n13771) );
  CMPR32X1 U21423 ( .A(n13772), .B(n13771), .C(n13770), .CO(n13834), .S(n13765) );
  ADDFHX1 U21424 ( .A(n13774), .B(n13775), .CI(n13773), .CO(n13853), .S(n13784) );
  OAI22XL U21425 ( .A0(n13776), .A1(n2997), .B0(n13899), .B1(n13844), .Y(
        n13847) );
  XNOR2XL U21426 ( .A(n14306), .B(n4807), .Y(n13840) );
  XNOR2XL U21427 ( .A(n4567), .B(n25863), .Y(n13837) );
  OAI22XL U21428 ( .A0(n13837), .A1(n14268), .B0(n13778), .B1(n14282), .Y(
        n13845) );
  XNOR2XL U21429 ( .A(n14288), .B(n14030), .Y(n13860) );
  OAI22XL U21430 ( .A0(n13860), .A1(n14029), .B0(n13779), .B1(n14044), .Y(
        n13859) );
  XNOR2XL U21431 ( .A(n14027), .B(n23173), .Y(n13836) );
  ADDFHX1 U21432 ( .A(n13784), .B(n13783), .CI(n13782), .CO(n13829), .S(n13763) );
  OAI21XL U21433 ( .A0(n13787), .A1(n13786), .B0(n13785), .Y(n13789) );
  NAND2X1 U21434 ( .A(n13789), .B(n13788), .Y(n13828) );
  XNOR2XL U21435 ( .A(n14235), .B(n14156), .Y(n13861) );
  XNOR2XL U21436 ( .A(n14265), .B(n25861), .Y(n13841) );
  OAI22XL U21437 ( .A0(n13841), .A1(n3173), .B0(n13793), .B1(n14080), .Y(
        n13848) );
  INVXL U21438 ( .A(n13810), .Y(n13808) );
  OAI2BB1X2 U21439 ( .A0N(n13811), .A1N(n13810), .B0(n13809), .Y(n13822) );
  ADDFHX4 U21440 ( .A(n13817), .B(n13816), .CI(n13815), .CO(n13983), .S(n13646) );
  ADDFHX4 U21441 ( .A(n13820), .B(n13819), .CI(n13818), .CO(n13987), .S(n13986) );
  XNOR2XL U21442 ( .A(n4565), .B(n23173), .Y(n13873) );
  OAI22XL U21443 ( .A0(n13836), .A1(n6191), .B0(n13873), .B1(n14298), .Y(
        n13891) );
  XNOR2XL U21444 ( .A(n14118), .B(M1_b_19_), .Y(n13900) );
  OAI22XL U21445 ( .A0(n13837), .A1(n14282), .B0(n13900), .B1(n14251), .Y(
        n13890) );
  XNOR2X1 U21446 ( .A(n14236), .B(n25862), .Y(n13875) );
  XNOR2XL U21447 ( .A(n14196), .B(n14228), .Y(n13901) );
  OAI22XL U21448 ( .A0(n13839), .A1(n14249), .B0(n13901), .B1(n14250), .Y(
        n13879) );
  XNOR2XL U21449 ( .A(n14357), .B(n4807), .Y(n13871) );
  OAI22XL U21450 ( .A0(n13840), .A1(n13971), .B0(n13871), .B1(n13972), .Y(
        n13878) );
  XNOR2XL U21451 ( .A(n25864), .B(n25861), .Y(n13874) );
  OAI22X1 U21452 ( .A0(n2993), .A1(n13919), .B0(n14289), .B1(n14028), .Y(
        n13896) );
  ADDFHX1 U21453 ( .A(n13847), .B(n13846), .CI(n13845), .CO(n13869), .S(n13852) );
  ADDFHX1 U21454 ( .A(n13859), .B(n13858), .CI(n13857), .CO(n13882), .S(n13851) );
  XNOR2XL U21455 ( .A(n14307), .B(n14030), .Y(n13872) );
  XNOR2XL U21456 ( .A(n14266), .B(n14156), .Y(n13876) );
  CMPR32X1 U21457 ( .A(n13864), .B(n13863), .C(n13862), .CO(n13892), .S(n13865) );
  CMPR32X1 U21458 ( .A(n13867), .B(n13866), .C(n13865), .CO(n13880), .S(n13835) );
  ADDFHX1 U21459 ( .A(n13870), .B(n13869), .CI(n13868), .CO(n13910), .S(n13886) );
  OAI22XL U21460 ( .A0(n13871), .A1(n13971), .B0(n13972), .B1(n4807), .Y(
        n13913) );
  OAI22X1 U21461 ( .A0(n13934), .A1(n14029), .B0(n13872), .B1(n14044), .Y(
        n13912) );
  XNOR2XL U21462 ( .A(n4567), .B(n23173), .Y(n13933) );
  OAI22XL U21463 ( .A0(n13933), .A1(n14291), .B0(n13873), .B1(n6191), .Y(
        n13911) );
  XNOR2XL U21464 ( .A(n14288), .B(n25861), .Y(n13932) );
  OAI22XL U21465 ( .A0(n13916), .A1(n14120), .B0(n13876), .B1(n14121), .Y(
        n13929) );
  CMPR32X1 U21466 ( .A(n13879), .B(n13878), .C(n13877), .CO(n13935), .S(n13887) );
  ADDFHX1 U21467 ( .A(n13882), .B(n13881), .CI(n13880), .CO(n13908), .S(n13902) );
  CMPR32X1 U21468 ( .A(n13888), .B(n13887), .C(n13886), .CO(n13940), .S(n13884) );
  CMPR32X1 U21469 ( .A(n13891), .B(n13890), .C(n13889), .CO(n13922), .S(n13888) );
  OAI22XL U21470 ( .A0(n2993), .A1(n14028), .B0(n14356), .B1(n14027), .Y(
        n13918) );
  XNOR2XL U21471 ( .A(n14195), .B(n14228), .Y(n13915) );
  OAI22X1 U21472 ( .A0(n13915), .A1(n14227), .B0(n13901), .B1(n14249), .Y(
        n13926) );
  ADDFHX1 U21473 ( .A(n13904), .B(n13903), .CI(n13902), .CO(n13938), .S(n13883) );
  ADDFHX1 U21474 ( .A(n13913), .B(n13912), .CI(n13911), .CO(n13955), .S(n13937) );
  XNOR2XL U21475 ( .A(n14266), .B(n25862), .Y(n13976) );
  XNOR2XL U21476 ( .A(n25864), .B(n14156), .Y(n13962) );
  CMPR32X1 U21477 ( .A(n25865), .B(n13919), .C(n13918), .CO(n13965), .S(n13925) );
  OAI22X1 U21478 ( .A0(n2993), .A1(n14027), .B0(n14356), .B1(n4565), .Y(n13968) );
  OAI22XL U21479 ( .A0(n13971), .A1(n4807), .B0(n13972), .B1(n13047), .Y(
        n13967) );
  XNOR2XL U21480 ( .A(n14307), .B(n25861), .Y(n13977) );
  OAI22XL U21481 ( .A0(n13932), .A1(n14080), .B0(n13977), .B1(n3173), .Y(
        n13958) );
  XNOR2XL U21482 ( .A(n14118), .B(n23173), .Y(n13970) );
  ADDFHX4 U21483 ( .A(n13943), .B(n13942), .CI(n13941), .CO(n13996), .S(n13995) );
  ADDFHX1 U21484 ( .A(n13949), .B(n13948), .CI(n13947), .CO(n14004), .S(n13950) );
  CMPR32X1 U21485 ( .A(n13955), .B(n13954), .C(n13953), .CO(n14010), .S(n13952) );
  XNOR2XL U21486 ( .A(n14288), .B(n14156), .Y(n14014) );
  XNOR2XL U21487 ( .A(n14235), .B(n14228), .Y(n14023) );
  CMPR32X1 U21488 ( .A(n13966), .B(n13965), .C(n13964), .CO(n14007), .S(n13953) );
  XNOR2XL U21489 ( .A(n14117), .B(n23173), .Y(n14024) );
  OAI22XL U21490 ( .A0(n14024), .A1(n14298), .B0(n13970), .B1(n6191), .Y(
        n14033) );
  OAI2BB1X1 U21491 ( .A0N(n13972), .A1N(n13971), .B0(n4807), .Y(n14032) );
  OAI22XL U21492 ( .A0(n14025), .A1(n14268), .B0(n13973), .B1(n14282), .Y(
        n14031) );
  XNOR2XL U21493 ( .A(n14306), .B(n25861), .Y(n14015) );
  OAI22XL U21494 ( .A0(n14015), .A1(n3173), .B0(n13977), .B1(n14080), .Y(
        n14011) );
  OAI21X2 U21495 ( .A0(n14618), .A1(n14632), .B0(n14619), .Y(n13991) );
  ADDFHX1 U21496 ( .A(n14004), .B(n14003), .CI(n14002), .CO(n14310), .S(n13998) );
  ADDFHX1 U21497 ( .A(n14007), .B(n14005), .CI(n14006), .CO(n14039), .S(n14008) );
  XNOR2XL U21498 ( .A(n14307), .B(n14156), .Y(n14058) );
  OAI22XL U21499 ( .A0(n14015), .A1(n14080), .B0(n14057), .B1(n3173), .Y(
        n14052) );
  CMPR32X1 U21500 ( .A(n14019), .B(n14018), .C(n14017), .CO(n14054), .S(n14020) );
  XNOR2XL U21501 ( .A(n14196), .B(n23173), .Y(n14047) );
  CMPR32X1 U21502 ( .A(n14028), .B(n14027), .C(n14026), .CO(n14065), .S(n14017) );
  ADDFHX1 U21503 ( .A(n14036), .B(n14035), .CI(n14034), .CO(n14040), .S(n14006) );
  OAI22XL U21504 ( .A0(n14075), .A1(n14198), .B0(n14046), .B1(n14208), .Y(
        n14094) );
  OAI22XL U21505 ( .A0(n14071), .A1(n14291), .B0(n14047), .B1(n6191), .Y(
        n14093) );
  CMPR32X1 U21506 ( .A(n14053), .B(n14052), .C(n14051), .CO(n14105), .S(n14055) );
  OAI22XL U21507 ( .A0(n14070), .A1(n14120), .B0(n14058), .B1(n14121), .Y(
        n14097) );
  XNOR2X1 U21508 ( .A(n14265), .B(n14228), .Y(n14076) );
  OAI22XL U21509 ( .A0(n14069), .A1(n14268), .B0(n14059), .B1(n14282), .Y(
        n14074) );
  OAI22XL U21510 ( .A0(n2993), .A1(n14118), .B0(n14356), .B1(n14117), .Y(
        n14077) );
  ADDFHX1 U21511 ( .A(n14062), .B(n14061), .CI(n14060), .CO(n14072), .S(n14064) );
  ADDFHX1 U21512 ( .A(n14065), .B(n14064), .CI(n14063), .CO(n14164), .S(n14041) );
  XNOR2XL U21513 ( .A(n14236), .B(n23173), .Y(n14078) );
  XNOR2X1 U21514 ( .A(n25864), .B(n14228), .Y(n14088) );
  OAI22XL U21515 ( .A0(n14076), .A1(n14249), .B0(n14088), .B1(n14227), .Y(
        n14086) );
  CMPR32X1 U21516 ( .A(n4565), .B(n4567), .C(n14077), .CO(n14085), .S(n14073)
         );
  OAI22XL U21517 ( .A0(n2993), .A1(n14196), .B0(n14289), .B1(n14195), .Y(
        n14116) );
  XNOR2XL U21518 ( .A(n14235), .B(n23173), .Y(n14133) );
  OAI22XL U21519 ( .A0(n14133), .A1(n14298), .B0(n14078), .B1(n6191), .Y(
        n14128) );
  XNOR2XL U21520 ( .A(n14265), .B(M1_b_19_), .Y(n14135) );
  XOR2X1 U21521 ( .A(n14125), .B(n14129), .Y(n14082) );
  XOR2X1 U21522 ( .A(n14128), .B(n14082), .Y(n14122) );
  CMPR32X1 U21523 ( .A(n14087), .B(n14086), .C(n14085), .CO(n14111), .S(n14102) );
  XNOR2XL U21524 ( .A(n14288), .B(n14228), .Y(n14115) );
  OAI22XL U21525 ( .A0(n14115), .A1(n14227), .B0(n14088), .B1(n14249), .Y(
        n14131) );
  OAI22XL U21526 ( .A0(n14134), .A1(n14198), .B0(n14089), .B1(n14208), .Y(
        n14130) );
  CMPR32X1 U21527 ( .A(n14095), .B(n14094), .C(n14093), .CO(n14100), .S(n14107) );
  ADDFHX1 U21528 ( .A(n14101), .B(n14100), .CI(n14099), .CO(n14112), .S(n14169) );
  CMPR32X1 U21529 ( .A(n14107), .B(n14106), .C(n14105), .CO(n14167), .S(n14172) );
  OAI21XL U21530 ( .A0(n14110), .A1(n14111), .B0(n14108), .Y(n14109) );
  CMPR32X1 U21531 ( .A(n14118), .B(n14117), .C(n14116), .CO(n14146), .S(n14124) );
  OAI22XL U21532 ( .A0(n14121), .A1(n14156), .B0(n14120), .B1(n14119), .Y(
        n14150) );
  CMPR32X1 U21533 ( .A(n14124), .B(n14123), .C(n14122), .CO(n14143), .S(n14114) );
  CMPR32X1 U21534 ( .A(n14132), .B(n14131), .C(n14130), .CO(n14140), .S(n14110) );
  XNOR2XL U21535 ( .A(n14266), .B(n23173), .Y(n14149) );
  OAI22XL U21536 ( .A0(n14133), .A1(n6191), .B0(n14149), .B1(n14298), .Y(
        n14155) );
  ADDFHX1 U21537 ( .A(n14141), .B(n14140), .CI(n14139), .CO(n14181), .S(n14142) );
  OAI22XL U21538 ( .A0(n14189), .A1(n14291), .B0(n14149), .B1(n6191), .Y(
        n14192) );
  OAI2BB1XL U21539 ( .A0N(n14120), .A1N(n14157), .B0(n14156), .Y(n14201) );
  XNOR2XL U21540 ( .A(n14288), .B(M1_b_19_), .Y(n14188) );
  OAI22XL U21541 ( .A0(n14188), .A1(n14268), .B0(n14158), .B1(n14282), .Y(
        n14200) );
  CMPR32X1 U21542 ( .A(n14166), .B(n14165), .C(n14164), .CO(n14175), .S(n14170) );
  ADDFHX1 U21543 ( .A(n14184), .B(n14183), .CI(n14182), .CO(n14204), .S(n14185) );
  OAI22XL U21544 ( .A0(n14189), .A1(n6191), .B0(n14209), .B1(n14298), .Y(
        n14212) );
  CMPR32X1 U21545 ( .A(n14193), .B(n14192), .C(n14191), .CO(n14219), .S(n14186) );
  CMPR32X1 U21546 ( .A(n14196), .B(n14195), .C(n14194), .CO(n14207), .S(n14191) );
  CMPR32X1 U21547 ( .A(n14201), .B(n14200), .C(n14199), .CO(n14205), .S(n14182) );
  CMPR32X1 U21548 ( .A(n14204), .B(n14203), .C(n14202), .CO(n14326), .S(n14323) );
  XNOR2XL U21549 ( .A(n14288), .B(n23173), .Y(n14232) );
  OAI22XL U21550 ( .A0(n14232), .A1(n14291), .B0(n14209), .B1(n6191), .Y(
        n14230) );
  CMPR32X1 U21551 ( .A(n14213), .B(n14212), .C(n14211), .CO(n14238), .S(n14220) );
  CMPR32X1 U21552 ( .A(n14217), .B(n14216), .C(n14215), .CO(n14224), .S(n14206) );
  CMPR32X1 U21553 ( .A(n14220), .B(n14219), .C(n14218), .CO(n14221), .S(n14202) );
  CMPR32X1 U21554 ( .A(n14223), .B(n14222), .C(n14221), .CO(n14328), .S(n14325) );
  CMPR32X1 U21555 ( .A(n14231), .B(n14230), .C(n14229), .CO(n14255), .S(n14239) );
  XNOR2XL U21556 ( .A(n14307), .B(n23173), .Y(n14253) );
  CMPR32X1 U21557 ( .A(n14236), .B(n14235), .C(n14234), .CO(n14243), .S(n14225) );
  CMPR32X1 U21558 ( .A(n14245), .B(n14244), .C(n14243), .CO(n14259), .S(n14254) );
  CMPR32X1 U21559 ( .A(n14248), .B(n14247), .C(n14246), .CO(n14270), .S(n14256) );
  OAI22X1 U21560 ( .A0(n14252), .A1(n14282), .B0(n14251), .B1(n25863), .Y(
        n14261) );
  XNOR2XL U21561 ( .A(n14306), .B(n23173), .Y(n14263) );
  CMPR32X1 U21562 ( .A(n14256), .B(n14255), .C(n14254), .CO(n14257), .S(n14241) );
  CMPR32X1 U21563 ( .A(n14259), .B(n14258), .C(n14257), .CO(n14332), .S(n14329) );
  XNOR2XL U21564 ( .A(n14357), .B(n23173), .Y(n14283) );
  CMPR32X1 U21565 ( .A(n14266), .B(n14265), .C(n14264), .CO(n14280), .S(n14271) );
  CMPR32X1 U21566 ( .A(n14275), .B(n14274), .C(n14273), .CO(n14339), .S(n14331) );
  CMPR32X1 U21567 ( .A(n14278), .B(n14277), .C(n14276), .CO(n14286), .S(n14279) );
  CMPR32X1 U21568 ( .A(n14281), .B(n14280), .C(n14279), .CO(n14285), .S(n14274) );
  CMPR32X1 U21569 ( .A(n14286), .B(n14285), .C(n14284), .CO(n14341), .S(n14338) );
  CMPR32X1 U21570 ( .A(n25864), .B(n14288), .C(n14287), .CO(n14297), .S(n14292) );
  CMPR32X1 U21571 ( .A(n14294), .B(n14293), .C(n14292), .CO(n14295), .S(n14284) );
  CMPR32X1 U21572 ( .A(n14297), .B(n14296), .C(n14295), .CO(n14343), .S(n14340) );
  CMPR32X1 U21573 ( .A(n14301), .B(n14300), .C(n14299), .CO(n14302), .S(n14296) );
  CMPR32X1 U21574 ( .A(n14304), .B(n14303), .C(n14302), .CO(n14348), .S(n14342) );
  CMPR32X1 U21575 ( .A(n14307), .B(n14306), .C(n14305), .CO(n14355), .S(n14303) );
  OR2X2 U21576 ( .A(n14348), .B(n14347), .Y(n14679) );
  NAND2XL U21577 ( .A(n14319), .B(n14320), .Y(n14525) );
  INVXL U21578 ( .A(n14525), .Y(n14321) );
  NAND2XL U21579 ( .A(n14326), .B(n14325), .Y(n14546) );
  NAND2XL U21580 ( .A(n14330), .B(n14329), .Y(n14490) );
  INVXL U21581 ( .A(n14490), .Y(n14494) );
  AOI21XL U21582 ( .A0(n14272), .A1(n14494), .B0(n14333), .Y(n14334) );
  OAI21XL U21583 ( .A0(n14335), .A1(n14538), .B0(n14334), .Y(n14336) );
  AOI21X2 U21584 ( .A0(n14534), .A1(n14337), .B0(n14336), .Y(n14502) );
  OAI21XL U21585 ( .A0(n14514), .A1(n14509), .B0(n14515), .Y(n14645) );
  CMPR32X1 U21586 ( .A(n14355), .B(n14354), .C(n14353), .CO(n14360), .S(n14347) );
  OAI21XL U21587 ( .A0(n14390), .A1(n14389), .B0(n14392), .Y(n14364) );
  OAI21XL U21588 ( .A0(M1_U4_U1_enc_tree_2__4__16_), .A1(
        M1_U3_U1_enc_tree_2__4__16_), .B0(n14364), .Y(n14370) );
  NAND2XL U21589 ( .A(n3152), .B(n14400), .Y(n14401) );
  XOR2X1 U21590 ( .A(n14402), .B(n14401), .Y(n14474) );
  OAI21XL U21591 ( .A0(n22472), .A1(n26142), .B0(n24022), .Y(n14406) );
  AOI2BB1X1 U21592 ( .A0N(n26286), .A1N(n3115), .B0(n14406), .Y(n14700) );
  OAI21XL U21593 ( .A0(n22472), .A1(n25936), .B0(n25216), .Y(n14409) );
  AOI21XL U21594 ( .A0(y11[26]), .A1(n14417), .B0(n25215), .Y(n14411) );
  OAI21XL U21595 ( .A0(n22472), .A1(n25937), .B0(n25213), .Y(n14412) );
  AOI21XL U21596 ( .A0(y11[28]), .A1(n14417), .B0(n25212), .Y(n14414) );
  OAI21XL U21597 ( .A0(n22472), .A1(n25935), .B0(n25210), .Y(n14415) );
  AOI21XL U21598 ( .A0(n14417), .A1(y11[30]), .B0(n24021), .Y(n14418) );
  OAI21XL U21599 ( .A0(n26303), .A1(n3115), .B0(n14418), .Y(n14703) );
  NOR2X1 U21600 ( .A(n14693), .B(n14703), .Y(n24028) );
  NOR4XL U21601 ( .A(y10[25]), .B(y10[29]), .C(y10[28]), .D(y10[30]), .Y(
        n14422) );
  NOR4XL U21602 ( .A(y10[26]), .B(y10[23]), .C(y10[22]), .D(y10[21]), .Y(
        n14421) );
  NOR4XL U21603 ( .A(y10[20]), .B(y10[19]), .C(y10[18]), .D(y10[17]), .Y(
        n14420) );
  NOR3XL U21604 ( .A(y10[0]), .B(y10[24]), .C(y10[27]), .Y(n14419) );
  NOR4XL U21605 ( .A(y10[16]), .B(y10[15]), .C(y10[14]), .D(y10[13]), .Y(
        n14426) );
  NOR4XL U21606 ( .A(y10[12]), .B(y10[11]), .C(y10[10]), .D(y10[9]), .Y(n14425) );
  NOR4XL U21607 ( .A(y10[8]), .B(y10[7]), .C(y10[6]), .D(y10[5]), .Y(n14424)
         );
  NOR4XL U21608 ( .A(y10[4]), .B(y10[3]), .C(y10[2]), .D(y10[1]), .Y(n14423)
         );
  OAI21X2 U21609 ( .A0(n14429), .A1(n14428), .B0(n14427), .Y(n14456) );
  NAND4X1 U21610 ( .A(n14456), .B(n14455), .C(n14454), .D(n14453), .Y(n14713)
         );
  CMPR32X1 U21611 ( .A(n14716), .B(n14458), .C(n14457), .CO(n14658), .S(n25774) );
  CMPR32X1 U21612 ( .A(n14712), .B(n14460), .C(n14459), .CO(n14467), .S(n24410) );
  CMPR32X1 U21613 ( .A(n14714), .B(n14462), .C(n14461), .CO(n14463), .S(n24083) );
  CMPR32X1 U21614 ( .A(n14710), .B(n14466), .C(n14465), .CO(n14457), .S(n24105) );
  CMPR32X1 U21615 ( .A(n14709), .B(n14468), .C(n14467), .CO(n14465), .S(n24280) );
  NAND4BXL U21616 ( .AN(n25774), .B(n14471), .C(n14470), .D(n14469), .Y(n14472) );
  INVXL U21617 ( .A(n14473), .Y(n14654) );
  NOR2XL U21618 ( .A(n14487), .B(n14532), .Y(n14493) );
  INVXL U21619 ( .A(n14493), .Y(n14489) );
  INVXL U21620 ( .A(n14538), .Y(n14485) );
  INVXL U21621 ( .A(n14496), .Y(n14488) );
  NAND2XL U21622 ( .A(n14493), .B(n14495), .Y(n14498) );
  NOR2X1 U21623 ( .A(n14503), .B(n14532), .Y(n14644) );
  INVXL U21624 ( .A(n14644), .Y(n14505) );
  INVXL U21625 ( .A(n14647), .Y(n14504) );
  NAND2XL U21626 ( .A(n14644), .B(n14511), .Y(n14513) );
  NOR2XL U21627 ( .A(n20688), .B(n4752), .Y(n14519) );
  INVXL U21628 ( .A(n14550), .Y(n14568) );
  NOR2XL U21629 ( .A(n14568), .B(n14521), .Y(n14559) );
  NAND2XL U21630 ( .A(n14559), .B(n14564), .Y(n14524) );
  NAND2XL U21631 ( .A(n5501), .B(n14535), .Y(n14537) );
  NAND2X1 U21632 ( .A(n14539), .B(n14538), .Y(n14540) );
  INVXL U21633 ( .A(n14541), .Y(n14542) );
  INVXL U21634 ( .A(n14545), .Y(n14547) );
  NAND2X1 U21635 ( .A(n14547), .B(n14546), .Y(n14548) );
  AOI21XL U21636 ( .A0(n14552), .A1(n14570), .B0(n14551), .Y(n14553) );
  INVXL U21637 ( .A(n14559), .Y(n14562) );
  INVXL U21638 ( .A(n14560), .Y(n14561) );
  INVX1 U21639 ( .A(n14687), .Y(n19092) );
  NOR2X1 U21640 ( .A(n19096), .B(n19092), .Y(n14578) );
  OAI21X1 U21641 ( .A0(n14677), .A1(n14568), .B0(n14567), .Y(n14572) );
  INVXL U21642 ( .A(n14573), .Y(n14575) );
  NAND2X1 U21643 ( .A(n14575), .B(n14574), .Y(n14576) );
  XNOR2X4 U21644 ( .A(n14577), .B(n14576), .Y(n14661) );
  INVXL U21645 ( .A(n14595), .Y(n14579) );
  NOR2XL U21646 ( .A(n14579), .B(n14598), .Y(n14582) );
  INVXL U21647 ( .A(n14624), .Y(n14604) );
  NAND2XL U21648 ( .A(n14582), .B(n14604), .Y(n14584) );
  INVX1 U21649 ( .A(n14623), .Y(n14606) );
  INVXL U21650 ( .A(n14594), .Y(n14580) );
  OAI21XL U21651 ( .A0(n14580), .A1(n14598), .B0(n14599), .Y(n14581) );
  AOI21XL U21652 ( .A0(n14606), .A1(n14582), .B0(n14581), .Y(n14583) );
  OAI21XL U21653 ( .A0(n14584), .A1(n14638), .B0(n14583), .Y(n14589) );
  NAND2XL U21654 ( .A(n14587), .B(n14586), .Y(n14588) );
  XNOR2X1 U21655 ( .A(n14589), .B(n14588), .Y(n20975) );
  NAND2XL U21656 ( .A(n14604), .B(n14595), .Y(n14597) );
  AOI21XL U21657 ( .A0(n14606), .A1(n14595), .B0(n14594), .Y(n14596) );
  OAI21XL U21658 ( .A0(n14597), .A1(n14638), .B0(n14596), .Y(n14602) );
  XNOR2X1 U21659 ( .A(n14602), .B(n14601), .Y(n20330) );
  NAND2XL U21660 ( .A(n14604), .B(n14626), .Y(n14608) );
  INVXL U21661 ( .A(n14614), .Y(n14633) );
  NAND2XL U21662 ( .A(n14629), .B(n14633), .Y(n14617) );
  INVXL U21663 ( .A(n14632), .Y(n14615) );
  NAND2XL U21664 ( .A(n14620), .B(n14619), .Y(n14621) );
  XNOR2X1 U21665 ( .A(n14622), .B(n14621), .Y(n20980) );
  INVXL U21666 ( .A(n14629), .Y(n14631) );
  NAND2XL U21667 ( .A(n14633), .B(n14632), .Y(n14634) );
  NAND2X1 U21668 ( .A(n14641), .B(n14640), .Y(n14642) );
  NAND2XL U21669 ( .A(n14644), .B(n14646), .Y(n14649) );
  OAI21X1 U21670 ( .A0(n14677), .A1(n14649), .B0(n14648), .Y(n14653) );
  XNOR2X1 U21671 ( .A(n14653), .B(n14652), .Y(n14682) );
  AOI21XL U21672 ( .A0(n14660), .A1(n24304), .B0(n24025), .Y(n14659) );
  NOR2X1 U21673 ( .A(n24025), .B(n14660), .Y(n24034) );
  NAND3X1 U21674 ( .A(n14661), .B(n20330), .C(n20975), .Y(n14667) );
  NAND4BX2 U21675 ( .AN(n14664), .B(n20982), .C(n20327), .D(n23589), .Y(n14665) );
  AND3X4 U21676 ( .A(n23706), .B(n14669), .C(n14668), .Y(n14670) );
  NAND2XL U21677 ( .A(n5501), .B(n14673), .Y(n14676) );
  AOI21XL U21678 ( .A0(n14674), .A1(n14673), .B0(n14672), .Y(n14675) );
  OAI21X1 U21679 ( .A0(n14696), .A1(n14695), .B0(n14694), .Y(n24036) );
  OAI21XL U21680 ( .A0(n14723), .A1(n14722), .B0(n14721), .Y(n22477) );
  NOR2XL U21681 ( .A(n14725), .B(n20688), .Y(n14726) );
  NOR2X1 U21682 ( .A(n14727), .B(n23709), .Y(n14728) );
  AOI22XL U21683 ( .A0(n19346), .A1(w2[72]), .B0(n3062), .B1(w1[104]), .Y(
        n14730) );
  OAI21XL U21684 ( .A0(n3063), .A1(n25972), .B0(n14730), .Y(n14996) );
  AOI22XL U21685 ( .A0(n19349), .A1(y12[8]), .B0(n3062), .B1(temp3[8]), .Y(
        n14731) );
  OAI21XL U21686 ( .A0(n14833), .A1(n26535), .B0(n14731), .Y(n14995) );
  NOR2XL U21687 ( .A(n15075), .B(n14995), .Y(n14734) );
  AOI22XL U21688 ( .A0(n19346), .A1(w2[73]), .B0(n19216), .B1(w1[105]), .Y(
        n14732) );
  OAI21XL U21689 ( .A0(n3063), .A1(n25971), .B0(n14732), .Y(n14998) );
  AOI22XL U21690 ( .A0(n19346), .A1(y12[9]), .B0(n19216), .B1(temp3[9]), .Y(
        n14733) );
  OAI21XL U21691 ( .A0(n14833), .A1(n26533), .B0(n14733), .Y(n14997) );
  NOR2XL U21692 ( .A(n15097), .B(n14997), .Y(n14795) );
  AOI22XL U21693 ( .A0(n19346), .A1(w2[75]), .B0(n3026), .B1(w1[107]), .Y(
        n14735) );
  OAI21XL U21694 ( .A0(n3063), .A1(n25969), .B0(n14735), .Y(n15006) );
  INVX1 U21695 ( .A(n15006), .Y(n15413) );
  AOI22XL U21696 ( .A0(n19346), .A1(y12[11]), .B0(n3062), .B1(temp3[11]), .Y(
        n14736) );
  OAI21XL U21697 ( .A0(n14833), .A1(n26531), .B0(n14736), .Y(n15005) );
  AOI22XL U21698 ( .A0(n19346), .A1(w2[74]), .B0(n3026), .B1(w1[106]), .Y(
        n14737) );
  OAI21XL U21699 ( .A0(n3063), .A1(n25970), .B0(n14737), .Y(n15002) );
  AOI22XL U21700 ( .A0(n19346), .A1(y12[10]), .B0(n3062), .B1(temp3[10]), .Y(
        n14738) );
  OAI21XL U21701 ( .A0(n14833), .A1(n26532), .B0(n14738), .Y(n15001) );
  NOR2XL U21702 ( .A(n15406), .B(n15001), .Y(n14739) );
  AOI22XL U21703 ( .A0(n19346), .A1(w2[76]), .B0(n19216), .B1(w1[108]), .Y(
        n14741) );
  OAI21XL U21704 ( .A0(n3063), .A1(n25968), .B0(n14741), .Y(n14981) );
  AOI22XL U21705 ( .A0(n19346), .A1(y12[12]), .B0(n3026), .B1(temp3[12]), .Y(
        n14742) );
  OAI21XL U21706 ( .A0(n3063), .A1(n26530), .B0(n14742), .Y(n14980) );
  AOI22XL U21707 ( .A0(n19346), .A1(w2[77]), .B0(n3026), .B1(w1[109]), .Y(
        n14743) );
  OAI21XL U21708 ( .A0(n3063), .A1(n25967), .B0(n14743), .Y(n14983) );
  INVX1 U21709 ( .A(n14983), .Y(n15430) );
  AOI22XL U21710 ( .A0(n19346), .A1(y12[13]), .B0(n3062), .B1(temp3[13]), .Y(
        n14744) );
  OAI21XL U21711 ( .A0(n14833), .A1(n26529), .B0(n14744), .Y(n14982) );
  AOI22XL U21712 ( .A0(n19346), .A1(w2[79]), .B0(n19216), .B1(w1[111]), .Y(
        n14746) );
  OAI21XL U21713 ( .A0(n3063), .A1(n25965), .B0(n14746), .Y(n14989) );
  AOI22XL U21714 ( .A0(n19346), .A1(y12[15]), .B0(n3026), .B1(temp3[15]), .Y(
        n14747) );
  OAI21XL U21715 ( .A0(n3063), .A1(n26527), .B0(n14747), .Y(n14988) );
  INVX1 U21716 ( .A(n14987), .Y(n15435) );
  AOI22XL U21717 ( .A0(n19346), .A1(y12[14]), .B0(n3026), .B1(temp3[14]), .Y(
        n14748) );
  OAI21XL U21718 ( .A0(n14833), .A1(n26528), .B0(n14748), .Y(n14986) );
  AOI22XL U21719 ( .A0(n3027), .A1(w2[67]), .B0(n19161), .B1(w1[99]), .Y(
        n14752) );
  OAI21XL U21720 ( .A0(n19237), .A1(n25977), .B0(n14752), .Y(n15175) );
  AOI22XL U21721 ( .A0(n19346), .A1(y12[3]), .B0(n19161), .B1(temp3[3]), .Y(
        n14753) );
  OAI21XL U21722 ( .A0(n14833), .A1(n26541), .B0(n14753), .Y(n15174) );
  NOR2XL U21723 ( .A(n15206), .B(n15174), .Y(n14766) );
  AOI22XL U21724 ( .A0(n19346), .A1(w2[66]), .B0(n19161), .B1(w1[98]), .Y(
        n14754) );
  OAI21XL U21725 ( .A0(n19237), .A1(n25978), .B0(n14754), .Y(n15172) );
  AOI22XL U21726 ( .A0(n19346), .A1(y12[2]), .B0(n19161), .B1(temp3[2]), .Y(
        n14755) );
  OAI21XL U21727 ( .A0(n19237), .A1(n26542), .B0(n14755), .Y(n15171) );
  NOR2XL U21728 ( .A(n15191), .B(n15171), .Y(n14756) );
  NOR2XL U21729 ( .A(n14766), .B(n14756), .Y(n14769) );
  AOI22XL U21730 ( .A0(n3027), .A1(w2[65]), .B0(n19161), .B1(w1[97]), .Y(
        n14757) );
  OAI21XL U21731 ( .A0(n19237), .A1(n25979), .B0(n14757), .Y(n15228) );
  AOI22XL U21732 ( .A0(n3027), .A1(y12[1]), .B0(n19161), .B1(temp3[1]), .Y(
        n14758) );
  OAI21XL U21733 ( .A0(n19237), .A1(n26543), .B0(n14758), .Y(n15227) );
  NOR2XL U21734 ( .A(n15259), .B(n15227), .Y(n14763) );
  AOI22XL U21735 ( .A0(n3027), .A1(w2[64]), .B0(n19161), .B1(w1[96]), .Y(
        n14759) );
  OAI21XL U21736 ( .A0(n19237), .A1(n25980), .B0(n14759), .Y(n15226) );
  AOI22XL U21737 ( .A0(n3027), .A1(y12[0]), .B0(n19161), .B1(temp3[0]), .Y(
        n14760) );
  OAI21XL U21738 ( .A0(n19237), .A1(n26544), .B0(n14760), .Y(n15225) );
  NAND2XL U21739 ( .A(n15242), .B(n15225), .Y(n14762) );
  NAND2XL U21740 ( .A(n15259), .B(n15227), .Y(n14761) );
  OAI21XL U21741 ( .A0(n14763), .A1(n14762), .B0(n14761), .Y(n14768) );
  NAND2XL U21742 ( .A(n15191), .B(n15171), .Y(n14765) );
  NAND2XL U21743 ( .A(n15206), .B(n15174), .Y(n14764) );
  OAI21XL U21744 ( .A0(n14766), .A1(n14765), .B0(n14764), .Y(n14767) );
  AOI22XL U21745 ( .A0(n3027), .A1(w2[68]), .B0(n19161), .B1(w1[100]), .Y(
        n14770) );
  OAI21XL U21746 ( .A0(n3063), .A1(n25976), .B0(n14770), .Y(n15177) );
  AOI22XL U21747 ( .A0(n19346), .A1(y12[4]), .B0(n19161), .B1(temp3[4]), .Y(
        n14771) );
  OAI21XL U21748 ( .A0(n3063), .A1(n26540), .B0(n14771), .Y(n15176) );
  NOR2XL U21749 ( .A(n15222), .B(n15176), .Y(n14774) );
  AOI22XL U21750 ( .A0(n3027), .A1(w2[69]), .B0(n19161), .B1(w1[101]), .Y(
        n14772) );
  OAI21XL U21751 ( .A0(n3063), .A1(n25975), .B0(n14772), .Y(n15155) );
  AOI22XL U21752 ( .A0(n19346), .A1(y12[5]), .B0(n19161), .B1(temp3[5]), .Y(
        n14773) );
  OAI21XL U21753 ( .A0(n14833), .A1(n26539), .B0(n14773), .Y(n15154) );
  NOR2XL U21754 ( .A(n14774), .B(n14783), .Y(n14780) );
  AOI22XL U21755 ( .A0(n19346), .A1(w2[70]), .B0(n19161), .B1(w1[102]), .Y(
        n14775) );
  OAI21XL U21756 ( .A0(n3063), .A1(n25974), .B0(n14775), .Y(n15103) );
  AOI22XL U21757 ( .A0(n19235), .A1(y12[6]), .B0(n19161), .B1(temp3[6]), .Y(
        n14776) );
  OAI21XL U21758 ( .A0(n14833), .A1(n26538), .B0(n14776), .Y(n15102) );
  NOR2XL U21759 ( .A(n15126), .B(n15102), .Y(n14779) );
  AOI22XL U21760 ( .A0(n19346), .A1(w2[71]), .B0(n19216), .B1(w1[103]), .Y(
        n14777) );
  OAI21XL U21761 ( .A0(n14833), .A1(n25973), .B0(n14777), .Y(n15106) );
  AOI22XL U21762 ( .A0(n19346), .A1(y12[7]), .B0(n3026), .B1(temp3[7]), .Y(
        n14778) );
  OAI21XL U21763 ( .A0(n14833), .A1(n26537), .B0(n14778), .Y(n15105) );
  NAND2XL U21764 ( .A(n14780), .B(n14789), .Y(n14791) );
  NAND2XL U21765 ( .A(n15222), .B(n15176), .Y(n14782) );
  NAND2XL U21766 ( .A(n15169), .B(n15154), .Y(n14781) );
  OAI21XL U21767 ( .A0(n14783), .A1(n14782), .B0(n14781), .Y(n14788) );
  NAND2XL U21768 ( .A(n15126), .B(n15102), .Y(n14785) );
  NAND2XL U21769 ( .A(n15150), .B(n15105), .Y(n14784) );
  OAI21XL U21770 ( .A0(n14786), .A1(n14785), .B0(n14784), .Y(n14787) );
  NAND2XL U21771 ( .A(n15075), .B(n14995), .Y(n14794) );
  NAND2XL U21772 ( .A(n15097), .B(n14997), .Y(n14793) );
  OAI21XL U21773 ( .A0(n14795), .A1(n14794), .B0(n14793), .Y(n14800) );
  NAND2XL U21774 ( .A(n15406), .B(n15001), .Y(n14797) );
  NAND2XL U21775 ( .A(n15413), .B(n15005), .Y(n14796) );
  OAI21XL U21776 ( .A0(n14798), .A1(n14797), .B0(n14796), .Y(n14799) );
  AOI21XL U21777 ( .A0(n14801), .A1(n14800), .B0(n14799), .Y(n14813) );
  NAND2XL U21778 ( .A(n15422), .B(n14980), .Y(n14803) );
  NAND2XL U21779 ( .A(n15430), .B(n14982), .Y(n14802) );
  OAI21XL U21780 ( .A0(n14804), .A1(n14803), .B0(n14802), .Y(n14809) );
  NAND2XL U21781 ( .A(n15435), .B(n14986), .Y(n14806) );
  NAND2XL U21782 ( .A(n15440), .B(n14988), .Y(n14805) );
  OAI21XL U21783 ( .A0(n14807), .A1(n14806), .B0(n14805), .Y(n14808) );
  AOI21XL U21784 ( .A0(n14810), .A1(n14809), .B0(n14808), .Y(n14811) );
  AOI21X1 U21785 ( .A0(n14816), .A1(n14815), .B0(n14814), .Y(n14907) );
  AOI22XL U21786 ( .A0(n19346), .A1(w2[80]), .B0(n19216), .B1(w1[112]), .Y(
        n14817) );
  OAI21XL U21787 ( .A0(n3063), .A1(n25964), .B0(n14817), .Y(n15057) );
  AOI22XL U21788 ( .A0(n19346), .A1(y12[16]), .B0(n3026), .B1(temp3[16]), .Y(
        n14818) );
  OAI21XL U21789 ( .A0(n3063), .A1(n26526), .B0(n14818), .Y(n15056) );
  AOI22XL U21790 ( .A0(n19346), .A1(w2[81]), .B0(n3062), .B1(w1[113]), .Y(
        n14819) );
  OAI21XL U21791 ( .A0(n3063), .A1(n25963), .B0(n14819), .Y(n15059) );
  AOI22XL U21792 ( .A0(n19346), .A1(y12[17]), .B0(n3026), .B1(temp3[17]), .Y(
        n14820) );
  OAI21XL U21793 ( .A0(n3063), .A1(n26525), .B0(n14820), .Y(n15058) );
  AOI22XL U21794 ( .A0(n3027), .A1(w2[83]), .B0(n19216), .B1(w1[115]), .Y(
        n14822) );
  OAI21XL U21795 ( .A0(n3063), .A1(n25961), .B0(n14822), .Y(n15066) );
  AOI22XL U21796 ( .A0(n3027), .A1(y12[19]), .B0(n3026), .B1(temp3[19]), .Y(
        n14823) );
  OAI21XL U21797 ( .A0(n3063), .A1(n26523), .B0(n14823), .Y(n15065) );
  AOI22XL U21798 ( .A0(n19346), .A1(w2[82]), .B0(n3026), .B1(w1[114]), .Y(
        n14824) );
  OAI21XL U21799 ( .A0(n3063), .A1(n25962), .B0(n14824), .Y(n15063) );
  AOI22XL U21800 ( .A0(n19346), .A1(y12[18]), .B0(n3062), .B1(temp3[18]), .Y(
        n14825) );
  OAI21XL U21801 ( .A0(n3063), .A1(n26524), .B0(n14825), .Y(n15062) );
  AOI22XL U21802 ( .A0(n3027), .A1(w2[84]), .B0(n19216), .B1(w1[116]), .Y(
        n14828) );
  OAI21XL U21803 ( .A0(n3063), .A1(n25960), .B0(n14828), .Y(n15048) );
  AOI22XL U21804 ( .A0(n3027), .A1(y12[20]), .B0(n3062), .B1(temp3[20]), .Y(
        n14829) );
  OAI21XL U21805 ( .A0(n3063), .A1(n26522), .B0(n14829), .Y(n15047) );
  AOI22XL U21806 ( .A0(n19346), .A1(w2[85]), .B0(n3026), .B1(w1[117]), .Y(
        n14830) );
  OAI21XL U21807 ( .A0(n3063), .A1(n25959), .B0(n14830), .Y(n15050) );
  AOI22XL U21808 ( .A0(n3027), .A1(y12[21]), .B0(n3026), .B1(temp3[21]), .Y(
        n14831) );
  OAI21XL U21809 ( .A0(n3063), .A1(n26521), .B0(n14831), .Y(n15049) );
  OAI21XL U21810 ( .A0(n19237), .A1(n26192), .B0(n14834), .Y(n14947) );
  AOI22XL U21811 ( .A0(n3027), .A1(w2[86]), .B0(n19216), .B1(w1[118]), .Y(
        n14836) );
  OAI21XL U21812 ( .A0(n3063), .A1(n25958), .B0(n14836), .Y(n15053) );
  AOI22XL U21813 ( .A0(n19346), .A1(y12[22]), .B0(n3026), .B1(temp3[22]), .Y(
        n14837) );
  OAI21XL U21814 ( .A0(n3063), .A1(n26520), .B0(n14837), .Y(n15052) );
  NOR2X1 U21815 ( .A(n14878), .B(n14838), .Y(n14881) );
  AOI22XL U21816 ( .A0(w2[88]), .A1(n19349), .B0(n19216), .B1(w1[120]), .Y(
        n14841) );
  OAI21XL U21817 ( .A0(n19237), .A1(n26193), .B0(n14841), .Y(n14943) );
  AOI22XL U21818 ( .A0(y12[24]), .A1(n19349), .B0(n3026), .B1(temp3[24]), .Y(
        n14842) );
  OAI21XL U21819 ( .A0(n19237), .A1(n26501), .B0(n14842), .Y(n14942) );
  NOR2XL U21820 ( .A(n14919), .B(n14942), .Y(n14845) );
  AOI22XL U21821 ( .A0(w2[89]), .A1(n19346), .B0(n3062), .B1(w1[121]), .Y(
        n14843) );
  INVX1 U21822 ( .A(n14951), .Y(n14917) );
  AOI22XL U21823 ( .A0(w2[91]), .A1(n19346), .B0(n19161), .B1(w1[123]), .Y(
        n14846) );
  AOI22XL U21824 ( .A0(y12[27]), .A1(n3027), .B0(n19161), .B1(temp3[27]), .Y(
        n14847) );
  AOI22XL U21825 ( .A0(w2[90]), .A1(n19346), .B0(n3062), .B1(w1[122]), .Y(
        n14848) );
  OAI21XL U21826 ( .A0(n14833), .A1(n26194), .B0(n14848), .Y(n14955) );
  AOI22XL U21827 ( .A0(y12[26]), .A1(n3027), .B0(n19161), .B1(temp3[26]), .Y(
        n14849) );
  NOR2XL U21828 ( .A(n14915), .B(n14954), .Y(n14850) );
  AOI22XL U21829 ( .A0(w2[92]), .A1(n19349), .B0(n19216), .B1(w1[124]), .Y(
        n14852) );
  OAI21XL U21830 ( .A0(n19237), .A1(n26191), .B0(n14852), .Y(n14931) );
  INVX1 U21831 ( .A(n14931), .Y(n14911) );
  AOI22XL U21832 ( .A0(y12[28]), .A1(n19349), .B0(n3026), .B1(temp3[28]), .Y(
        n14853) );
  OAI21XL U21833 ( .A0(n19237), .A1(n26498), .B0(n14853), .Y(n14930) );
  OAI21XL U21834 ( .A0(n19237), .A1(n26188), .B0(n14854), .Y(n14935) );
  INVX1 U21835 ( .A(n14935), .Y(n14909) );
  OAI21XL U21836 ( .A0(n19237), .A1(n26499), .B0(n14855), .Y(n14934) );
  NAND2XL U21837 ( .A(n15461), .B(n15056), .Y(n14864) );
  NAND2XL U21838 ( .A(n15521), .B(n15058), .Y(n14863) );
  OAI21XL U21839 ( .A0(n14865), .A1(n14864), .B0(n14863), .Y(n14870) );
  NAND2XL U21840 ( .A(n15537), .B(n15062), .Y(n14867) );
  NAND2XL U21841 ( .A(n15542), .B(n15065), .Y(n14866) );
  OAI21XL U21842 ( .A0(n14868), .A1(n14867), .B0(n14866), .Y(n14869) );
  AOI21XL U21843 ( .A0(n14871), .A1(n14870), .B0(n14869), .Y(n14884) );
  NAND2XL U21844 ( .A(n15547), .B(n15047), .Y(n14873) );
  NAND2XL U21845 ( .A(n15552), .B(n15049), .Y(n14872) );
  OAI21XL U21846 ( .A0(n14874), .A1(n14873), .B0(n14872), .Y(n14880) );
  NAND2XL U21847 ( .A(n15557), .B(n15052), .Y(n14877) );
  NAND2XL U21848 ( .A(n14875), .B(n14946), .Y(n14876) );
  OAI21XL U21849 ( .A0(n14878), .A1(n14877), .B0(n14876), .Y(n14879) );
  AOI21XL U21850 ( .A0(n14881), .A1(n14880), .B0(n14879), .Y(n14882) );
  OAI21XL U21851 ( .A0(n14884), .A1(n14883), .B0(n14882), .Y(n14904) );
  NAND2XL U21852 ( .A(n14919), .B(n14942), .Y(n14886) );
  NAND2XL U21853 ( .A(n14917), .B(n14950), .Y(n14885) );
  OAI21XL U21854 ( .A0(n14887), .A1(n14886), .B0(n14885), .Y(n14892) );
  NAND2XL U21855 ( .A(n14915), .B(n14954), .Y(n14889) );
  NAND2XL U21856 ( .A(n14913), .B(n14926), .Y(n14888) );
  OAI21XL U21857 ( .A0(n14890), .A1(n14889), .B0(n14888), .Y(n14891) );
  AOI21XL U21858 ( .A0(n14893), .A1(n14892), .B0(n14891), .Y(n14901) );
  NAND2XL U21859 ( .A(n14911), .B(n14930), .Y(n14895) );
  NAND2XL U21860 ( .A(n14909), .B(n14934), .Y(n14894) );
  OAI21XL U21861 ( .A0(n14896), .A1(n14895), .B0(n14894), .Y(n14898) );
  INVX8 U21862 ( .A(n3101), .Y(n15558) );
  OAI21X2 U21863 ( .A0(n15558), .A1(n14909), .B0(n14908), .Y(n24431) );
  NAND2XL U21864 ( .A(n15190), .B(n14930), .Y(n14910) );
  OAI21XL U21865 ( .A0(n15558), .A1(n14911), .B0(n14910), .Y(n24401) );
  NAND2XL U21866 ( .A(n15190), .B(n14926), .Y(n14912) );
  OAI21XL U21867 ( .A0(n15558), .A1(n14913), .B0(n14912), .Y(n24293) );
  NAND2X1 U21868 ( .A(n15190), .B(n14946), .Y(n14920) );
  CMPR22X1 U21869 ( .A(n4793), .B(n14921), .CO(n15735), .S(n24399) );
  CMPR22X1 U21870 ( .A(n4791), .B(n14922), .CO(n14921), .S(n24291) );
  NAND2X1 U21871 ( .A(n14941), .B(n14923), .Y(n24020) );
  NAND2XL U21872 ( .A(n15190), .B(n14927), .Y(n14928) );
  OAI21XL U21873 ( .A0(n15558), .A1(n14933), .B0(n14932), .Y(n23159) );
  OAI21XL U21874 ( .A0(n15558), .A1(n14941), .B0(n14940), .Y(n23157) );
  NAND2XL U21875 ( .A(n15190), .B(n14955), .Y(n14956) );
  NOR2X1 U21876 ( .A(n24100), .B(n14968), .Y(n14974) );
  OAI21X2 U21877 ( .A0(n14974), .A1(n14977), .B0(n14975), .Y(n15015) );
  NOR2X1 U21878 ( .A(n24355), .B(n14969), .Y(n15010) );
  NOR2X1 U21879 ( .A(n4787), .B(n14970), .Y(n15013) );
  INVXL U21880 ( .A(n15013), .Y(n14971) );
  INVXL U21881 ( .A(n14974), .Y(n14976) );
  NAND2XL U21882 ( .A(n14976), .B(n14975), .Y(n14978) );
  XOR2X1 U21883 ( .A(n14978), .B(n14977), .Y(n15128) );
  XNOR2X1 U21884 ( .A(n23966), .B(n14979), .Y(n15004) );
  NAND2XL U21885 ( .A(n3038), .B(n14984), .Y(n14985) );
  OAI21XL U21886 ( .A0(n3038), .A1(n15338), .B0(n14985), .Y(n15099) );
  OAI21XL U21887 ( .A0(n15008), .A1(n15441), .B0(n14990), .Y(n15324) );
  NAND2XL U21888 ( .A(n3038), .B(n15324), .Y(n14991) );
  OAI21XL U21889 ( .A0(n3038), .A1(n15302), .B0(n14991), .Y(n15118) );
  NAND2XL U21890 ( .A(n15055), .B(n14992), .Y(n14993) );
  OAI21XL U21891 ( .A0(n15055), .A1(n15099), .B0(n14993), .Y(n15209) );
  INVXL U21892 ( .A(n15010), .Y(n14994) );
  NAND2XL U21893 ( .A(n3038), .B(n14999), .Y(n15000) );
  OAI21XL U21894 ( .A0(n3038), .A1(n15288), .B0(n15000), .Y(n15108) );
  OAI21XL U21895 ( .A0(n15558), .A1(n15407), .B0(n15003), .Y(n15279) );
  OAI21XL U21896 ( .A0(n15008), .A1(n15414), .B0(n15007), .Y(n15323) );
  AOI22XL U21897 ( .A0(n15289), .A1(n15279), .B0(n3038), .B1(n15323), .Y(
        n15101) );
  NAND2XL U21898 ( .A(n15055), .B(n15101), .Y(n15009) );
  OAI21XL U21899 ( .A0(n15055), .A1(n15108), .B0(n15009), .Y(n15213) );
  OAI22XL U21900 ( .A0(n15209), .A1(n6194), .B0(n3016), .B1(n15213), .Y(n15236) );
  NOR2XL U21901 ( .A(n15010), .B(n15013), .Y(n15016) );
  OAI21XL U21902 ( .A0(n15045), .A1(n15041), .B0(n15042), .Y(n15021) );
  NAND2XL U21903 ( .A(n4793), .B(n15018), .Y(n15022) );
  OAI21XL U21904 ( .A0(n15023), .A1(n15042), .B0(n15022), .Y(n15035) );
  INVXL U21905 ( .A(n15035), .Y(n15025) );
  NOR2XL U21906 ( .A(n15023), .B(n15041), .Y(n15032) );
  INVXL U21907 ( .A(n15032), .Y(n15024) );
  NAND2XL U21908 ( .A(n15032), .B(n15026), .Y(n15037) );
  AOI21XL U21909 ( .A0(n15035), .A1(n15026), .B0(n15034), .Y(n15036) );
  OAI21XL U21910 ( .A0(n15045), .A1(n15037), .B0(n15036), .Y(n15039) );
  INVXL U21911 ( .A(n15041), .Y(n15043) );
  XOR2X2 U21912 ( .A(n15045), .B(n15044), .Y(n15355) );
  OAI21XL U21913 ( .A0(n15558), .A1(n15553), .B0(n15051), .Y(n15317) );
  AOI22XL U21914 ( .A0(n15289), .A1(n15089), .B0(n3038), .B1(n15317), .Y(
        n15112) );
  OAI21XL U21915 ( .A0(n15558), .A1(n15559), .B0(n15054), .Y(n15315) );
  OAI21XL U21916 ( .A0(n15558), .A1(n15522), .B0(n15060), .Y(n15275) );
  NAND2XL U21917 ( .A(n3038), .B(n15275), .Y(n15061) );
  OAI21XL U21918 ( .A0(n3038), .A1(n15334), .B0(n15061), .Y(n15115) );
  OAI21XL U21919 ( .A0(n15558), .A1(n15538), .B0(n15064), .Y(n15314) );
  OAI21XL U21920 ( .A0(n15558), .A1(n15543), .B0(n15067), .Y(n15283) );
  NAND2XL U21921 ( .A(n3038), .B(n15283), .Y(n15068) );
  OAI21XL U21922 ( .A0(n3038), .A1(n15069), .B0(n15068), .Y(n15114) );
  INVXL U21923 ( .A(n15114), .Y(n15070) );
  NAND2XL U21924 ( .A(n15055), .B(n15070), .Y(n15071) );
  OAI21XL U21925 ( .A0(n15055), .A1(n15115), .B0(n15071), .Y(n15210) );
  INVX1 U21926 ( .A(n23955), .Y(n15364) );
  AOI21XL U21927 ( .A0(n15074), .A1(n23955), .B0(n15573), .Y(n15073) );
  NAND2XL U21928 ( .A(n3038), .B(n15077), .Y(n15078) );
  OAI21XL U21929 ( .A0(n3038), .A1(n15320), .B0(n15078), .Y(n15135) );
  AOI22XL U21930 ( .A0(n15289), .A1(n15324), .B0(n3038), .B1(n15079), .Y(
        n15131) );
  NAND2XL U21931 ( .A(n15055), .B(n15131), .Y(n15080) );
  OAI21XL U21932 ( .A0(n15055), .A1(n15135), .B0(n15080), .Y(n15152) );
  OAI21XL U21933 ( .A0(n3038), .A1(n15304), .B0(n15081), .Y(n15142) );
  NAND2XL U21934 ( .A(n15004), .B(n15082), .Y(n15083) );
  OAI21XL U21935 ( .A0(n3038), .A1(n15084), .B0(n15083), .Y(n15138) );
  INVXL U21936 ( .A(n15138), .Y(n15085) );
  NAND2XL U21937 ( .A(n15055), .B(n15085), .Y(n15086) );
  OAI21XL U21938 ( .A0(n15055), .A1(n15142), .B0(n15086), .Y(n15159) );
  OAI22XL U21939 ( .A0(n15152), .A1(n3156), .B0(n3016), .B1(n15159), .Y(n15252) );
  AOI22XL U21940 ( .A0(n15289), .A1(n15317), .B0(n3038), .B1(n15315), .Y(
        n15132) );
  NAND2XL U21941 ( .A(n3038), .B(n15314), .Y(n15087) );
  OAI21XL U21942 ( .A0(n3038), .A1(n15088), .B0(n15087), .Y(n15129) );
  NAND2XL U21943 ( .A(n3038), .B(n15089), .Y(n15090) );
  OAI21XL U21944 ( .A0(n3038), .A1(n15091), .B0(n15090), .Y(n15134) );
  INVXL U21945 ( .A(n15134), .Y(n15092) );
  NAND2XL U21946 ( .A(n15055), .B(n15092), .Y(n15093) );
  OAI21XL U21947 ( .A0(n15055), .A1(n15129), .B0(n15093), .Y(n15153) );
  AOI21XL U21948 ( .A0(n15096), .A1(n23955), .B0(n15573), .Y(n15095) );
  OAI21XL U21949 ( .A0(n14967), .A1(n15096), .B0(n15095), .Y(n15396) );
  INVXL U21950 ( .A(n15099), .Y(n15100) );
  AOI22XL U21951 ( .A0(n3167), .A1(n15101), .B0(n15100), .B1(n15055), .Y(
        n15182) );
  OAI21XL U21952 ( .A0(n15558), .A1(n15127), .B0(n15104), .Y(n15301) );
  OAI21XL U21953 ( .A0(n15558), .A1(n15151), .B0(n15107), .Y(n15290) );
  AOI22XL U21954 ( .A0(n15289), .A1(n15301), .B0(n3038), .B1(n15290), .Y(
        n15211) );
  INVXL U21955 ( .A(n15211), .Y(n15111) );
  INVXL U21956 ( .A(n15108), .Y(n15109) );
  NAND2XL U21957 ( .A(n15055), .B(n15109), .Y(n15110) );
  OAI21XL U21958 ( .A0(n15055), .A1(n15111), .B0(n15110), .Y(n15179) );
  AOI2BB2XL U21959 ( .B0(n15182), .B1(n3016), .A0N(n3016), .A1N(n15179), .Y(
        n15268) );
  NAND2XL U21960 ( .A(n15055), .B(n15112), .Y(n15113) );
  OAI21XL U21961 ( .A0(n15055), .A1(n15114), .B0(n15113), .Y(n15183) );
  INVXL U21962 ( .A(n15183), .Y(n15119) );
  INVXL U21963 ( .A(n15115), .Y(n15116) );
  NAND2XL U21964 ( .A(n15055), .B(n15116), .Y(n15117) );
  OAI21XL U21965 ( .A0(n15055), .A1(n15118), .B0(n15117), .Y(n15181) );
  INVXL U21966 ( .A(n15129), .Y(n15130) );
  AOI22XL U21967 ( .A0(n3167), .A1(n15131), .B0(n15130), .B1(n15055), .Y(
        n15199) );
  NAND2XL U21968 ( .A(n15055), .B(n15132), .Y(n15133) );
  OAI21XL U21969 ( .A0(n15055), .A1(n15134), .B0(n15133), .Y(n15200) );
  INVXL U21970 ( .A(n15135), .Y(n15136) );
  NAND2XL U21971 ( .A(n15055), .B(n15136), .Y(n15137) );
  OAI21XL U21972 ( .A0(n15055), .A1(n15138), .B0(n15137), .Y(n15198) );
  INVXL U21973 ( .A(n15290), .Y(n15141) );
  NAND2XL U21974 ( .A(n3038), .B(n15139), .Y(n15140) );
  OAI21XL U21975 ( .A0(n3038), .A1(n15141), .B0(n15140), .Y(n15157) );
  NAND2XL U21976 ( .A(n15055), .B(n15143), .Y(n15144) );
  OAI21XL U21977 ( .A0(n15055), .A1(n15157), .B0(n15144), .Y(n15195) );
  CLKINVX2 U21978 ( .A(n15355), .Y(n15340) );
  OAI21XL U21979 ( .A0(n15358), .A1(n3090), .B0(n15340), .Y(n15145) );
  AOI21XL U21980 ( .A0(n15149), .A1(n23955), .B0(n15573), .Y(n15148) );
  NAND2XL U21981 ( .A(n15558), .B(n15155), .Y(n15156) );
  OAI21XL U21982 ( .A0(n15558), .A1(n15170), .B0(n15156), .Y(n15327) );
  AOI22XL U21983 ( .A0(n15289), .A1(n15327), .B0(n3038), .B1(n15301), .Y(
        n15194) );
  INVXL U21984 ( .A(n15157), .Y(n15158) );
  AOI22XL U21985 ( .A0(n3167), .A1(n15194), .B0(n15158), .B1(n15055), .Y(
        n15248) );
  OAI21XL U21986 ( .A0(n15427), .A1(n3034), .B0(n15163), .Y(n15164) );
  OAI21XL U21987 ( .A0(n15558), .A1(n15192), .B0(n15173), .Y(n15325) );
  AOI22XL U21988 ( .A0(n15289), .A1(n15325), .B0(n3038), .B1(n15193), .Y(
        n15231) );
  OAI21XL U21989 ( .A0(n15558), .A1(n15223), .B0(n15178), .Y(n15294) );
  AOI22XL U21990 ( .A0(n15289), .A1(n15294), .B0(n3038), .B1(n15327), .Y(
        n15212) );
  AOI22XL U21991 ( .A0(n3167), .A1(n15231), .B0(n15212), .B1(n15055), .Y(
        n15265) );
  AOI21XL U21992 ( .A0(n15180), .A1(n15313), .B0(n15355), .Y(n15186) );
  NAND2XL U21993 ( .A(n15402), .B(n3090), .Y(n15185) );
  NOR2X1 U21994 ( .A(n15401), .B(n3090), .Y(n15534) );
  AOI22XL U21995 ( .A0(n15186), .A1(n15185), .B0(n15534), .B1(n15355), .Y(
        n15187) );
  AOI21XL U21996 ( .A0(n15189), .A1(n23955), .B0(n15573), .Y(n15188) );
  OAI21XL U21997 ( .A0(n14967), .A1(n15189), .B0(n15188), .Y(n15374) );
  NOR2XL U21998 ( .A(n15374), .B(n15373), .Y(n15648) );
  INVXL U21999 ( .A(n15648), .Y(n15653) );
  AOI22XL U22000 ( .A0(n15289), .A1(n15193), .B0(n3038), .B1(n15294), .Y(
        n15246) );
  INVXL U22001 ( .A(n15195), .Y(n15196) );
  AOI22XL U22002 ( .A0(n15354), .A1(n6194), .B0(n15196), .B1(n3016), .Y(n15197) );
  AOI21XL U22003 ( .A0(n15197), .A1(n15313), .B0(n15355), .Y(n15202) );
  NAND2XL U22004 ( .A(n15409), .B(n3090), .Y(n15201) );
  NAND2XL U22005 ( .A(n3167), .B(n15289), .Y(n15277) );
  AOI2BB2X1 U22006 ( .B0(n15303), .B1(n3016), .A0N(n3016), .A1N(n15200), .Y(
        n15408) );
  AOI22XL U22007 ( .A0(n15202), .A1(n15201), .B0(n15539), .B1(n15355), .Y(
        n15203) );
  AOI21XL U22008 ( .A0(n15205), .A1(n23955), .B0(n15573), .Y(n15204) );
  OAI21XL U22009 ( .A0(n14967), .A1(n15205), .B0(n15204), .Y(n15376) );
  NAND2XL U22010 ( .A(n15653), .B(n15208), .Y(n15642) );
  AOI22XL U22011 ( .A0(n3167), .A1(n15212), .B0(n15211), .B1(n15055), .Y(
        n15232) );
  OAI21XL U22012 ( .A0(n15419), .A1(n3034), .B0(n15216), .Y(n15217) );
  NOR2XL U22013 ( .A(n15224), .B(n3090), .Y(n15458) );
  INVXL U22014 ( .A(n15458), .Y(n15238) );
  INVXL U22015 ( .A(n15305), .Y(n15230) );
  INVXL U22016 ( .A(n15306), .Y(n15229) );
  AOI22XL U22017 ( .A0(n3167), .A1(n15264), .B0(n15231), .B1(n15055), .Y(
        n15233) );
  AOI22XL U22018 ( .A0(n15233), .A1(n3156), .B0(n15232), .B1(n3016), .Y(n15234) );
  AOI21XL U22019 ( .A0(n15234), .A1(n3034), .B0(n15355), .Y(n15235) );
  OAI21XL U22020 ( .A0(n3034), .A1(n15236), .B0(n15235), .Y(n15237) );
  OAI21XL U22021 ( .A0(n15238), .A1(n15340), .B0(n15237), .Y(n15239) );
  NAND2XL U22022 ( .A(n15256), .B(n15239), .Y(n15241) );
  AOI21XL U22023 ( .A0(n15241), .A1(n23955), .B0(n15573), .Y(n15240) );
  OAI21XL U22024 ( .A0(n14967), .A1(n15241), .B0(n15240), .Y(n15367) );
  OR2X2 U22025 ( .A(n15367), .B(n15366), .Y(n15691) );
  INVXL U22026 ( .A(n15518), .Y(n15254) );
  NAND2XL U22027 ( .A(n15004), .B(n15325), .Y(n15245) );
  OAI21XL U22028 ( .A0(n3038), .A1(n15306), .B0(n15245), .Y(n15351) );
  AOI22XL U22029 ( .A0(n3167), .A1(n15247), .B0(n15246), .B1(n15055), .Y(
        n15249) );
  AOI22XL U22030 ( .A0(n15249), .A1(n6194), .B0(n15248), .B1(n3016), .Y(n15250) );
  AOI21XL U22031 ( .A0(n15250), .A1(n15313), .B0(n15355), .Y(n15251) );
  OAI21XL U22032 ( .A0(n3034), .A1(n15252), .B0(n15251), .Y(n15253) );
  OAI21XL U22033 ( .A0(n15254), .A1(n15340), .B0(n15253), .Y(n15255) );
  NAND2XL U22034 ( .A(n15256), .B(n15255), .Y(n15258) );
  AOI21XL U22035 ( .A0(n15258), .A1(n23955), .B0(n15573), .Y(n15257) );
  OAI21XL U22036 ( .A0(n14967), .A1(n15258), .B0(n15257), .Y(n15369) );
  NAND2XL U22037 ( .A(n15691), .B(n15261), .Y(n15372) );
  AOI22XL U22038 ( .A0(n15266), .A1(n6194), .B0(n15265), .B1(n3016), .Y(n15267) );
  AOI21XL U22039 ( .A0(n15267), .A1(n3034), .B0(n15355), .Y(n15270) );
  NAND2XL U22040 ( .A(n15268), .B(n3090), .Y(n15269) );
  AOI22XL U22041 ( .A0(n15355), .A1(n15432), .B0(n15270), .B1(n15269), .Y(
        n15271) );
  NOR2XL U22042 ( .A(n15271), .B(n15359), .Y(n15273) );
  NAND2XL U22043 ( .A(n15273), .B(n15415), .Y(n15272) );
  OAI211XL U22044 ( .A0(n15364), .A1(n15273), .B0(n15363), .C0(n15272), .Y(
        n15274) );
  INVXL U22045 ( .A(n15336), .Y(n15276) );
  AOI211XL U22046 ( .A0(n15276), .A1(n15275), .B0(n15325), .C0(n15301), .Y(
        n15287) );
  OAI21XL U22047 ( .A0(n3034), .A1(n15312), .B0(n15340), .Y(n15280) );
  AOI21XL U22048 ( .A0(n15280), .A1(n15279), .B0(n15278), .Y(n15286) );
  AOI21XL U22049 ( .A0(n3034), .A1(n15289), .B0(n15281), .Y(n15284) );
  AOI211XL U22050 ( .A0(n3034), .A1(n3167), .B0(n15336), .C0(n15340), .Y(
        n15282) );
  OAI21XL U22051 ( .A0(n15284), .A1(n15283), .B0(n15282), .Y(n15285) );
  OAI211XL U22052 ( .A0(n15340), .A1(n15287), .B0(n15286), .C0(n15285), .Y(
        n15300) );
  NOR2XL U22053 ( .A(n15355), .B(n3016), .Y(n15293) );
  AOI21XL U22054 ( .A0(n15293), .A1(n15289), .B0(n15288), .Y(n15291) );
  NOR2XL U22055 ( .A(n15291), .B(n15290), .Y(n15292) );
  NOR2XL U22056 ( .A(n15355), .B(n3090), .Y(n15307) );
  AOI211XL U22057 ( .A0(n15293), .A1(n3167), .B0(n15292), .C0(n15307), .Y(
        n15299) );
  INVXL U22058 ( .A(n15307), .Y(n15328) );
  OAI21XL U22059 ( .A0(n15328), .A1(n3038), .B0(n15294), .Y(n15297) );
  AOI22XL U22060 ( .A0(n15297), .A1(n15296), .B0(n15307), .B1(n15295), .Y(
        n15298) );
  NOR3XL U22061 ( .A(n15300), .B(n15299), .C(n15298), .Y(n15347) );
  AOI22XL U22062 ( .A0(n15316), .A1(n15301), .B0(n15352), .B1(n15055), .Y(
        n15311) );
  AOI211XL U22063 ( .A0(n15336), .A1(n15303), .B0(n15302), .C0(n15340), .Y(
        n15310) );
  NAND2XL U22064 ( .A(n3090), .B(n3016), .Y(n15322) );
  AOI21XL U22065 ( .A0(n15322), .A1(n15340), .B0(n15304), .Y(n15309) );
  AOI22XL U22066 ( .A0(n15307), .A1(n3156), .B0(n15306), .B1(n15305), .Y(
        n15308) );
  NAND2XL U22067 ( .A(n15313), .B(n15312), .Y(n15326) );
  AOI22XL U22068 ( .A0(n15316), .A1(n15315), .B0(n15326), .B1(n15314), .Y(
        n15321) );
  OAI21XL U22069 ( .A0(n15318), .A1(n15317), .B0(n3090), .Y(n15319) );
  AOI31XL U22070 ( .A0(n15321), .A1(n15320), .A2(n15319), .B0(n15340), .Y(
        n15332) );
  AOI21XL U22071 ( .A0(n15336), .A1(n3167), .B0(n15340), .Y(n15333) );
  OAI21XL U22072 ( .A0(n15322), .A1(n3167), .B0(n15340), .Y(n15337) );
  AOI22XL U22073 ( .A0(n15328), .A1(n15327), .B0(n15326), .B1(n15325), .Y(
        n15330) );
  NAND4BXL U22074 ( .AN(n15332), .B(n15331), .C(n15330), .D(n15329), .Y(n15343) );
  INVXL U22075 ( .A(n15333), .Y(n15335) );
  AOI211XL U22076 ( .A0(n15336), .A1(n15289), .B0(n15335), .C0(n15334), .Y(
        n15342) );
  INVXL U22077 ( .A(n15337), .Y(n15339) );
  AOI211XL U22078 ( .A0(n15340), .A1(n15289), .B0(n15339), .C0(n15338), .Y(
        n15341) );
  AOI22XL U22079 ( .A0(n15350), .A1(n3090), .B0(n15349), .B1(n15313), .Y(
        n15437) );
  NAND2XL U22080 ( .A(n15437), .B(n15355), .Y(n15361) );
  AOI22XL U22081 ( .A0(n3167), .A1(n15352), .B0(n15055), .B1(n15351), .Y(
        n15353) );
  AOI21XL U22082 ( .A0(n15356), .A1(n15313), .B0(n15355), .Y(n15357) );
  OAI21XL U22083 ( .A0(n3034), .A1(n15358), .B0(n15357), .Y(n15360) );
  AOI21XL U22084 ( .A0(n15361), .A1(n15360), .B0(n15359), .Y(n15365) );
  NAND2XL U22085 ( .A(n15365), .B(n15415), .Y(n15362) );
  OAI211XL U22086 ( .A0(n15365), .A1(n15364), .B0(n15363), .C0(n15362), .Y(
        n15694) );
  NAND2XL U22087 ( .A(n15367), .B(n15366), .Y(n15690) );
  INVXL U22088 ( .A(n15690), .Y(n15657) );
  NAND2XL U22089 ( .A(n15369), .B(n15368), .Y(n15658) );
  INVXL U22090 ( .A(n15658), .Y(n15370) );
  INVXL U22091 ( .A(n15652), .Y(n15378) );
  NAND2XL U22092 ( .A(n15376), .B(n15375), .Y(n15649) );
  INVXL U22093 ( .A(n15649), .Y(n15377) );
  OAI21XL U22094 ( .A0(n15641), .A1(n15643), .B0(n15644), .Y(n15381) );
  OAI21XL U22095 ( .A0(n15512), .A1(n15670), .B0(n15513), .Y(n15397) );
  AOI21XL U22096 ( .A0(n15405), .A1(n23955), .B0(n15573), .Y(n15404) );
  OAI21XL U22097 ( .A0(n14967), .A1(n15405), .B0(n15404), .Y(n15443) );
  AOI21XL U22098 ( .A0(n15412), .A1(n23955), .B0(n15573), .Y(n15411) );
  OAI21XL U22099 ( .A0(n14967), .A1(n15412), .B0(n15411), .Y(n15445) );
  OAI21XL U22100 ( .A0(n15417), .A1(n3016), .B0(n3090), .Y(n15418) );
  AOI21XL U22101 ( .A0(n15421), .A1(n23955), .B0(n15573), .Y(n15420) );
  OAI21XL U22102 ( .A0(n14967), .A1(n15421), .B0(n15420), .Y(n15447) );
  OAI21XL U22103 ( .A0(n15425), .A1(n3016), .B0(n3090), .Y(n15426) );
  AOI21XL U22104 ( .A0(n15429), .A1(n23955), .B0(n15573), .Y(n15428) );
  OAI21XL U22105 ( .A0(n14967), .A1(n15429), .B0(n15428), .Y(n15449) );
  AOI21XL U22106 ( .A0(n15434), .A1(n23955), .B0(n15573), .Y(n15433) );
  OAI21XL U22107 ( .A0(n14967), .A1(n15434), .B0(n15433), .Y(n15453) );
  AOI21XL U22108 ( .A0(n15439), .A1(n23955), .B0(n15573), .Y(n15438) );
  OAI21XL U22109 ( .A0(n14967), .A1(n15439), .B0(n15438), .Y(n15455) );
  OAI21XL U22110 ( .A0(n15498), .A1(n15504), .B0(n15499), .Y(n15491) );
  OAI21XL U22111 ( .A0(n15485), .A1(n15494), .B0(n15486), .Y(n15450) );
  OAI21XL U22112 ( .A0(n15472), .A1(n15477), .B0(n15473), .Y(n15604) );
  AOI21XL U22113 ( .A0(n15610), .A1(n15601), .B0(n15604), .Y(n15456) );
  OAI21XL U22114 ( .A0(n15613), .A1(n15457), .B0(n15456), .Y(n15467) );
  AOI21XL U22115 ( .A0(n15460), .A1(n23955), .B0(n15573), .Y(n15459) );
  OAI21XL U22116 ( .A0(n14967), .A1(n15460), .B0(n15459), .Y(n15464) );
  NOR2X1 U22117 ( .A(n15464), .B(n15463), .Y(n15606) );
  OAI21XL U22118 ( .A0(n15613), .A1(n15471), .B0(n15470), .Y(n15476) );
  OAI21XL U22119 ( .A0(n15613), .A1(n15523), .B0(n15530), .Y(n15480) );
  AOI21XL U22120 ( .A0(n15491), .A1(n15495), .B0(n15482), .Y(n15483) );
  OAI21XL U22121 ( .A0(n15613), .A1(n15484), .B0(n15483), .Y(n15489) );
  OAI21XL U22122 ( .A0(n15613), .A1(n15493), .B0(n15492), .Y(n15497) );
  OAI21XL U22123 ( .A0(n15613), .A1(n15503), .B0(n15504), .Y(n15502) );
  OAI21XL U22124 ( .A0(n15509), .A1(n15669), .B0(n15670), .Y(n15510) );
  AOI21XL U22125 ( .A0(n15520), .A1(n23955), .B0(n15573), .Y(n15519) );
  OAI21XL U22126 ( .A0(n15614), .A1(n15605), .B0(n15615), .Y(n15526) );
  OAI21XL U22127 ( .A0(n14967), .A1(n15536), .B0(n15535), .Y(n15561) );
  AOI21XL U22128 ( .A0(n15541), .A1(n23955), .B0(n15573), .Y(n15540) );
  AOI21XL U22129 ( .A0(n15546), .A1(n23955), .B0(n15573), .Y(n15545) );
  AOI21XL U22130 ( .A0(n15551), .A1(n23955), .B0(n15573), .Y(n15550) );
  OR2X2 U22131 ( .A(n15620), .B(n15580), .Y(n15584) );
  OAI21XL U22132 ( .A0(n15633), .A1(n15626), .B0(n15634), .Y(n15568) );
  AOI21XL U22133 ( .A0(n15575), .A1(n23955), .B0(n15573), .Y(n15574) );
  OAI21XL U22134 ( .A0(n15619), .A1(n15580), .B0(n15576), .Y(n15577) );
  OAI21XL U22135 ( .A0(n15632), .A1(n15588), .B0(n15587), .Y(n15591) );
  OAI21XL U22136 ( .A0(n15632), .A1(n15597), .B0(n15598), .Y(n15596) );
  OAI21XL U22137 ( .A0(n15607), .A1(n15606), .B0(n15605), .Y(n15608) );
  OAI21XL U22138 ( .A0(n15613), .A1(n15612), .B0(n15611), .Y(n15618) );
  OAI21XL U22139 ( .A0(n15632), .A1(n15620), .B0(n15619), .Y(n15624) );
  AOI21XL U22140 ( .A0(n15629), .A1(n15628), .B0(n15627), .Y(n15630) );
  OAI21XL U22141 ( .A0(n15632), .A1(n15631), .B0(n15630), .Y(n15637) );
  CMPR22X1 U22142 ( .A(n4787), .B(n15639), .CO(n14922), .S(n24058) );
  OAI21XL U22143 ( .A0(n15655), .A1(n15642), .B0(n15641), .Y(n15647) );
  XNOR2X1 U22144 ( .A(n15651), .B(n15650), .Y(n15823) );
  XOR2X1 U22145 ( .A(n15655), .B(n15654), .Y(n15835) );
  INVXL U22146 ( .A(n15656), .Y(n15693) );
  AOI21XL U22147 ( .A0(n15693), .A1(n15691), .B0(n15657), .Y(n15660) );
  NAND2XL U22148 ( .A(n15261), .B(n15658), .Y(n15659) );
  XOR2X1 U22149 ( .A(n15660), .B(n15659), .Y(n15836) );
  AOI21XL U22150 ( .A0(n15680), .A1(n15665), .B0(n15661), .Y(n15664) );
  XOR2X1 U22151 ( .A(n15664), .B(n15663), .Y(n15819) );
  AOI21XL U22152 ( .A0(n15680), .A1(n15668), .B0(n15667), .Y(n15673) );
  OAI21XL U22153 ( .A0(n15677), .A1(n15676), .B0(n15675), .Y(n15678) );
  AOI21XL U22154 ( .A0(n15680), .A1(n15679), .B0(n15678), .Y(n15684) );
  CMPR22X1 U22155 ( .A(n24355), .B(n15689), .CO(n15639), .S(n24353) );
  NAND2XL U22156 ( .A(n15691), .B(n15690), .Y(n15692) );
  INVXL U22157 ( .A(n15694), .Y(n15696) );
  XNOR2XL U22158 ( .A(n15696), .B(n15695), .Y(n15754) );
  OAI21XL U22159 ( .A0(n15699), .A1(n15698), .B0(n15697), .Y(n15701) );
  INVXL U22160 ( .A(n15772), .Y(n15705) );
  AOI2BB1XL U22161 ( .A0N(n15820), .A1N(n15707), .B0(n15819), .Y(n15708) );
  AOI2BB1XL U22162 ( .A0N(n15708), .A1N(n15809), .B0(n15801), .Y(n15709) );
  INVXL U22163 ( .A(n15709), .Y(n15711) );
  INVXL U22164 ( .A(n15827), .Y(n15710) );
  AOI21XL U22165 ( .A0(n15711), .A1(n15710), .B0(n15826), .Y(n15712) );
  INVXL U22166 ( .A(n15873), .Y(n15713) );
  INVXL U22167 ( .A(n15715), .Y(n15717) );
  INVXL U22168 ( .A(n24870), .Y(n15716) );
  OAI21XL U22169 ( .A0(n15772), .A1(n15754), .B0(n15718), .Y(n15719) );
  OAI21XL U22170 ( .A0(n15723), .A1(n15722), .B0(n15721), .Y(n15724) );
  CMPR22X1 U22171 ( .A(n24100), .B(n23966), .CO(n15689), .S(n24098) );
  NOR3X1 U22172 ( .A(n24426), .B(n24399), .C(n15742), .Y(n15739) );
  CMPR22X1 U22173 ( .A(n24431), .B(n15735), .CO(n15736), .S(n24426) );
  CMPR22X1 U22174 ( .A(n24020), .B(n15736), .CO(n15737), .S(n24018) );
  XOR2X1 U22175 ( .A(n24426), .B(n15740), .Y(n24429) );
  CMPR32X1 U22176 ( .A(n24353), .B(n15745), .C(n15744), .CO(n15743), .S(n24354) );
  ADDFHX1 U22177 ( .A(n15746), .B(n25273), .CI(n24098), .CO(n15744), .S(n24099) );
  NOR4XL U22178 ( .A(n24059), .B(n24354), .C(n23964), .D(n24099), .Y(n15749)
         );
  INVXL U22179 ( .A(n24292), .Y(n15748) );
  OAI21XL U22180 ( .A0(n25269), .A1(n15753), .B0(n15752), .Y(n15807) );
  OAI21XL U22181 ( .A0(n25269), .A1(n23956), .B0(n15756), .Y(n15760) );
  NAND2XL U22182 ( .A(n15760), .B(n25273), .Y(n15853) );
  NOR2XL U22183 ( .A(n15853), .B(n24917), .Y(n15890) );
  NAND4BXL U22184 ( .AN(n15771), .B(n25007), .C(n24870), .D(n24962), .Y(n15780) );
  INVXL U22185 ( .A(n24020), .Y(n15788) );
  INVXL U22186 ( .A(n24431), .Y(n15787) );
  NAND4XL U22187 ( .A(n4792), .B(n15788), .C(n15787), .D(n23965), .Y(n15791)
         );
  NOR2XL U22188 ( .A(n24100), .B(n24355), .Y(n15789) );
  NAND3XL U22189 ( .A(n15789), .B(n4786), .C(n4790), .Y(n15790) );
  NAND4XL U22190 ( .A(n15818), .B(n15794), .C(n15793), .D(n15792), .Y(n15795)
         );
  NOR2X2 U22191 ( .A(n23963), .B(n15795), .Y(n24617) );
  NAND2XL U22192 ( .A(n25271), .B(n15872), .Y(n15796) );
  OAI21XL U22193 ( .A0(n25269), .A1(n15797), .B0(n15796), .Y(n15912) );
  NAND2XL U22194 ( .A(n25271), .B(n15860), .Y(n15798) );
  OAI21XL U22195 ( .A0(n25269), .A1(n15713), .B0(n15798), .Y(n15884) );
  OAI22XL U22196 ( .A0(n3127), .A1(n15912), .B0(n15884), .B1(n3070), .Y(n24874) );
  NAND2XL U22197 ( .A(n25271), .B(n15826), .Y(n15799) );
  OAI21XL U22198 ( .A0(n25269), .A1(n15800), .B0(n15799), .Y(n15883) );
  NOR2XL U22199 ( .A(n25269), .B(n15710), .Y(n15803) );
  NAND2XL U22200 ( .A(n15843), .B(n3127), .Y(n15804) );
  OAI21XL U22201 ( .A0(n3127), .A1(n15883), .B0(n15804), .Y(n15852) );
  OAI22XL U22202 ( .A0(n15808), .A1(n24874), .B0(n15852), .B1(n3125), .Y(
        n25265) );
  NOR2XL U22203 ( .A(n25265), .B(n15688), .Y(n15817) );
  OAI21XL U22204 ( .A0(n25271), .A1(n15806), .B0(n15805), .Y(n15848) );
  OAI22XL U22205 ( .A0(n3127), .A1(n15848), .B0(n15807), .B1(n3070), .Y(n15854) );
  NAND2XL U22206 ( .A(n25271), .B(n15819), .Y(n15810) );
  OAI21XL U22207 ( .A0(n25269), .A1(n15831), .B0(n15810), .Y(n15845) );
  NOR2XL U22208 ( .A(n25271), .B(n15811), .Y(n15813) );
  NAND2XL U22209 ( .A(n15846), .B(n3127), .Y(n15814) );
  OAI21XL U22210 ( .A0(n3127), .A1(n15845), .B0(n15814), .Y(n15851) );
  NOR2XL U22211 ( .A(n15891), .B(n3077), .Y(n15816) );
  NAND2XL U22212 ( .A(n25271), .B(n15820), .Y(n15821) );
  OAI21XL U22213 ( .A0(n25271), .A1(n15822), .B0(n15821), .Y(n15865) );
  NAND2XL U22214 ( .A(n25271), .B(n15823), .Y(n15824) );
  OAI21XL U22215 ( .A0(n25269), .A1(n15825), .B0(n15824), .Y(n15857) );
  OAI22XL U22216 ( .A0(n3127), .A1(n15865), .B0(n15857), .B1(n3070), .Y(n15878) );
  OAI21XL U22217 ( .A0(n25271), .A1(n15829), .B0(n15828), .Y(n15864) );
  NOR2XL U22218 ( .A(n25271), .B(n15830), .Y(n15833) );
  NAND2XL U22219 ( .A(n15866), .B(n3127), .Y(n15834) );
  OAI21XL U22220 ( .A0(n3127), .A1(n15864), .B0(n15834), .Y(n15876) );
  OAI22XL U22221 ( .A0(n15878), .A1(n3125), .B0(n15876), .B1(n15808), .Y(
        n21008) );
  NAND2XL U22222 ( .A(n25271), .B(n15836), .Y(n15837) );
  OAI21XL U22223 ( .A0(n25271), .A1(n15838), .B0(n15837), .Y(n15856) );
  NAND2XL U22224 ( .A(n15839), .B(n3127), .Y(n15840) );
  OAI21XL U22225 ( .A0(n3127), .A1(n15856), .B0(n15840), .Y(n15877) );
  NOR2XL U22226 ( .A(n15900), .B(n3077), .Y(n15841) );
  NAND2XL U22227 ( .A(n15843), .B(n25273), .Y(n15844) );
  OAI21XL U22228 ( .A0(n15845), .A1(n3070), .B0(n15844), .Y(n15885) );
  NAND2XL U22229 ( .A(n15846), .B(n25273), .Y(n15847) );
  OAI21XL U22230 ( .A0(n15848), .A1(n3070), .B0(n15847), .Y(n15881) );
  OAI22XL U22231 ( .A0(n15808), .A1(n15885), .B0(n15881), .B1(n3125), .Y(
        n15909) );
  OAI22XL U22232 ( .A0(n15808), .A1(n15852), .B0(n15851), .B1(n15745), .Y(
        n24869) );
  OAI22XL U22233 ( .A0(n15854), .A1(n15808), .B0(n3125), .B1(n15853), .Y(
        n15898) );
  OAI22XL U22234 ( .A0(n3127), .A1(n15857), .B0(n15856), .B1(n3070), .Y(n15892) );
  NAND2XL U22235 ( .A(n15858), .B(n24917), .Y(n15859) );
  OAI21XL U22236 ( .A0(n15892), .A1(n15808), .B0(n15859), .Y(n15899) );
  NAND2XL U22237 ( .A(n25271), .B(n15861), .Y(n15862) );
  OAI21XL U22238 ( .A0(n25269), .A1(n15863), .B0(n15862), .Y(n15875) );
  OAI22XL U22239 ( .A0(n3127), .A1(n15875), .B0(n15864), .B1(n3070), .Y(n15927) );
  INVXL U22240 ( .A(n15865), .Y(n15867) );
  AOI22XL U22241 ( .A0(n15867), .A1(n3127), .B0(n15866), .B1(n3070), .Y(n15893) );
  NAND2XL U22242 ( .A(n15893), .B(n24917), .Y(n15868) );
  OAI21XL U22243 ( .A0(n15808), .A1(n15927), .B0(n15868), .Y(n24925) );
  NOR2XL U22244 ( .A(n24925), .B(n15688), .Y(n15869) );
  NAND2XL U22245 ( .A(n24637), .B(n24663), .Y(n15871) );
  INVXL U22246 ( .A(n24667), .Y(n24773) );
  NAND2XL U22247 ( .A(n25271), .B(n15873), .Y(n15874) );
  OAI21XL U22248 ( .A0(n25269), .A1(n3138), .B0(n15874), .Y(n15924) );
  OAI22XL U22249 ( .A0(n3127), .A1(n15924), .B0(n15875), .B1(n25273), .Y(
        n21005) );
  OAI22XL U22250 ( .A0(n15808), .A1(n21005), .B0(n15876), .B1(n3125), .Y(
        n25006) );
  OAI22XL U22251 ( .A0(n15808), .A1(n15878), .B0(n15877), .B1(n3125), .Y(
        n15888) );
  NOR2XL U22252 ( .A(n15888), .B(n3077), .Y(n15879) );
  OAI22XL U22253 ( .A0(n3125), .A1(n15882), .B0(n15881), .B1(n15808), .Y(
        n15889) );
  NOR2XL U22254 ( .A(n15889), .B(n3077), .Y(n15887) );
  OAI22XL U22255 ( .A0(n3127), .A1(n15884), .B0(n15883), .B1(n3070), .Y(n15913) );
  OAI22XL U22256 ( .A0(n15808), .A1(n15913), .B0(n15885), .B1(n15745), .Y(
        n24971) );
  NOR2XL U22257 ( .A(n24971), .B(n15688), .Y(n15886) );
  NAND2XL U22258 ( .A(n24703), .B(n24670), .Y(n24770) );
  NOR2XL U22259 ( .A(n24773), .B(n24770), .Y(n15903) );
  NOR2XL U22260 ( .A(n25019), .B(n15638), .Y(n24541) );
  NAND2XL U22261 ( .A(n15889), .B(n3077), .Y(n24973) );
  NOR2XL U22262 ( .A(n24973), .B(n15638), .Y(n24518) );
  NAND2XL U22263 ( .A(n15894), .B(n15688), .Y(n15895) );
  NAND2XL U22264 ( .A(n15895), .B(n3076), .Y(n15896) );
  NAND2XL U22265 ( .A(n24584), .B(n24591), .Y(n15897) );
  NAND2XL U22266 ( .A(n15898), .B(n3077), .Y(n24877) );
  NAND2XL U22267 ( .A(n15899), .B(n3077), .Y(n24927) );
  NOR2XL U22268 ( .A(n24927), .B(n15638), .Y(n24507) );
  NAND2XL U22269 ( .A(n24502), .B(n24507), .Y(n15901) );
  NOR2XL U22270 ( .A(n21009), .B(n15638), .Y(n24469) );
  NAND2XL U22271 ( .A(n24469), .B(n25138), .Y(n24482) );
  NAND2XL U22272 ( .A(n15903), .B(n24775), .Y(n15905) );
  XOR2X1 U22273 ( .A(n15905), .B(n15904), .Y(n15906) );
  OAI21XL U22274 ( .A0(n25059), .A1(n25931), .B0(n15907), .Y(n15908) );
  AOI2BB1XL U22275 ( .A0N(n25461), .A1N(n3118), .B0(n15908), .Y(n2214) );
  NOR2XL U22276 ( .A(n15909), .B(n3077), .Y(n15918) );
  NAND2XL U22277 ( .A(n25271), .B(n15920), .Y(n15910) );
  OAI21XL U22278 ( .A0(n25269), .A1(n15911), .B0(n15910), .Y(n24873) );
  OAI22XL U22279 ( .A0(n3127), .A1(n24873), .B0(n15912), .B1(n3070), .Y(n24967) );
  OAI21XL U22280 ( .A0(n24967), .A1(n15808), .B0(n3077), .Y(n15915) );
  NOR2XL U22281 ( .A(n15913), .B(n3125), .Y(n15914) );
  OAI22XL U22282 ( .A0(n15918), .A1(n15917), .B0(n15916), .B1(n3076), .Y(
        n24881) );
  INVXL U22283 ( .A(n15919), .Y(n15932) );
  NOR2XL U22284 ( .A(n25269), .B(n15921), .Y(n15922) );
  AOI21XL U22285 ( .A0(n15923), .A1(n25269), .B0(n15922), .Y(n21003) );
  NOR2XL U22286 ( .A(n15924), .B(n3070), .Y(n15925) );
  AOI21XL U22287 ( .A0(n21003), .A1(n3070), .B0(n15925), .Y(n24914) );
  NAND2XL U22288 ( .A(n3125), .B(n24914), .Y(n15926) );
  OAI21XL U22289 ( .A0(n3125), .A1(n15927), .B0(n15926), .Y(n15930) );
  NAND2XL U22290 ( .A(n15928), .B(n15688), .Y(n15929) );
  OAI21XL U22291 ( .A0(n3076), .A1(n15932), .B0(n15931), .Y(n24780) );
  NAND2XL U22292 ( .A(n24771), .B(n24780), .Y(n15933) );
  NOR2XL U22293 ( .A(n15933), .B(n24770), .Y(n15934) );
  NOR2X2 U22294 ( .A(n15936), .B(n15935), .Y(n25286) );
  XNOR2XL U22295 ( .A(n25286), .B(n4781), .Y(n15937) );
  AOI22X1 U22296 ( .A0(n3029), .A1(n4782), .B0(n25290), .B1(n15937), .Y(n25437) );
  OAI21XL U22297 ( .A0(n25059), .A1(n26274), .B0(n15938), .Y(n15939) );
  AOI2BB1XL U22298 ( .A0N(n25437), .A1N(n3118), .B0(n15939), .Y(n2216) );
  OAI222X2 U22299 ( .A0(n26038), .A1(n15942), .B0(n26280), .B1(n25767), .C0(
        n25923), .C1(n15940), .Y(M5_a_20_) );
  XNOR2X1 U22300 ( .A(n3211), .B(n16884), .Y(n15955) );
  OAI22XL U22301 ( .A0(n16701), .A1(n15998), .B0(n16699), .B1(n15958), .Y(
        n15990) );
  NAND2X1 U22302 ( .A(n15948), .B(n16332), .Y(n16330) );
  XNOR2X1 U22303 ( .A(n16289), .B(n3201), .Y(n15964) );
  XNOR2X1 U22304 ( .A(n16289), .B(n3196), .Y(n15959) );
  XNOR2XL U22305 ( .A(n3203), .B(n12701), .Y(n15983) );
  OAI22XL U22306 ( .A0(n16867), .A1(n15973), .B0(n16939), .B1(n15983), .Y(
        n15987) );
  XOR2X1 U22307 ( .A(M5_a_12_), .B(n3199), .Y(n15950) );
  NAND2X2 U22308 ( .A(n15950), .B(n15996), .Y(n16893) );
  XNOR2XL U22309 ( .A(n3199), .B(M3_mult_x_15_b_13_), .Y(n15961) );
  OAI22X1 U22310 ( .A0(n16977), .A1(n16001), .B0(n3105), .B1(n15961), .Y(
        n15953) );
  XNOR2XL U22311 ( .A(n3022), .B(n11499), .Y(n16003) );
  XNOR2X1 U22312 ( .A(n3022), .B(n2974), .Y(n15962) );
  ADDFHX1 U22313 ( .A(n15953), .B(n15952), .CI(n3205), .CO(n16149), .S(n16041)
         );
  XNOR2X1 U22314 ( .A(n17039), .B(M3_mult_x_15_b_9_), .Y(n15960) );
  OAI22X1 U22315 ( .A0(n17060), .A1(n15960), .B0(n17061), .B1(n16127), .Y(
        n16133) );
  XNOR2X1 U22316 ( .A(n3211), .B(n3190), .Y(n15954) );
  XNOR2X1 U22317 ( .A(n3203), .B(n3198), .Y(n15982) );
  XNOR2XL U22318 ( .A(n3203), .B(n11495), .Y(n16142) );
  OAI22XL U22319 ( .A0(n16867), .A1(n15982), .B0(n16939), .B1(n16142), .Y(
        n16131) );
  XNOR2XL U22320 ( .A(n16614), .B(M3_mult_x_15_b_21_), .Y(n15957) );
  INVX8 U22321 ( .A(n16605), .Y(n16614) );
  OAI22XL U22322 ( .A0(n16701), .A1(n15957), .B0(n16699), .B1(n16125), .Y(
        n16129) );
  OAI22XL U22323 ( .A0(n16701), .A1(n15958), .B0(n16699), .B1(n15957), .Y(
        n16032) );
  XNOR2X1 U22324 ( .A(n17073), .B(M3_mult_x_15_b_6_), .Y(n16005) );
  XNOR2XL U22325 ( .A(n5677), .B(n3197), .Y(n15963) );
  OAI22XL U22326 ( .A0(n17074), .A1(n16005), .B0(n16375), .B1(n15963), .Y(
        n16030) );
  XNOR2X1 U22327 ( .A(n3022), .B(M3_mult_x_15_b_6_), .Y(n16135) );
  OAI22X1 U22328 ( .A0(n17092), .A1(n15962), .B0(n16317), .B1(n16135), .Y(
        n16122) );
  OAI22XL U22329 ( .A0(n17074), .A1(n15963), .B0(n16375), .B1(n16128), .Y(
        n16121) );
  XNOR2XL U22330 ( .A(n16289), .B(n11495), .Y(n16009) );
  XNOR2X1 U22331 ( .A(n17039), .B(M3_mult_x_15_b_6_), .Y(n16008) );
  OAI22XL U22332 ( .A0(n17060), .A1(n16008), .B0(n17061), .B1(n15966), .Y(
        n16052) );
  XNOR2XL U22333 ( .A(n15968), .B(n11495), .Y(n15979) );
  OAI22XL U22334 ( .A0(n17148), .A1(M3_mult_x_15_b_1_), .B0(n17147), .B1(
        M3_mult_x_15_b_2_), .Y(n15981) );
  NOR2BX1 U22335 ( .AN(n3110), .B(n17147), .Y(n16016) );
  OAI22X2 U22336 ( .A0(n16686), .A1(n16012), .B0(n15971), .B1(n16475), .Y(
        n16015) );
  XNOR2X1 U22337 ( .A(n3022), .B(M3_mult_x_15_b_1_), .Y(n16064) );
  OAI22X1 U22338 ( .A0(n16686), .A1(n15971), .B0(n16475), .B1(M5_mult_x_15_n1), 
        .Y(n15986) );
  XNOR2X1 U22339 ( .A(n3022), .B(M3_mult_x_15_b_3_), .Y(n16004) );
  XNOR2X1 U22340 ( .A(n17073), .B(n2974), .Y(n16006) );
  OAI22XL U22341 ( .A0(n17074), .A1(n16007), .B0(n16375), .B1(n16006), .Y(
        n15984) );
  XNOR2XL U22342 ( .A(n15968), .B(n12701), .Y(n16011) );
  XNOR2X1 U22343 ( .A(n3203), .B(n12561), .Y(n16010) );
  CMPR22X1 U22344 ( .A(n15975), .B(n15974), .CO(n15977), .S(n15999) );
  XNOR2X1 U22345 ( .A(n15968), .B(n3201), .Y(n16020) );
  CMPR32X1 U22346 ( .A(n3110), .B(n15981), .C(n15980), .CO(n16024), .S(n15976)
         );
  OAI22XL U22347 ( .A0(n17148), .A1(M3_mult_x_15_b_2_), .B0(n17147), .B1(
        n12279), .Y(n16022) );
  OAI22XL U22348 ( .A0(n16941), .A1(n15983), .B0(n16939), .B1(n15982), .Y(
        n16021) );
  ADDFHX1 U22349 ( .A(n15986), .B(n15985), .CI(n15984), .CO(n15995), .S(n16061) );
  OAI22X1 U22350 ( .A0(n16977), .A1(n16047), .B0(n3105), .B1(n16002), .Y(
        n16056) );
  XNOR2X1 U22351 ( .A(n16614), .B(n3196), .Y(n16050) );
  OAI22XL U22352 ( .A0(n16701), .A1(n16050), .B0(n16699), .B1(n15998), .Y(
        n16054) );
  OAI22X1 U22353 ( .A0(n16977), .A1(n16002), .B0(n3105), .B1(n16001), .Y(
        n16028) );
  OAI22XL U22354 ( .A0(n17074), .A1(n16006), .B0(n16375), .B1(n16005), .Y(
        n16026) );
  XNOR2XL U22355 ( .A(n3211), .B(n3197), .Y(n16069) );
  XNOR2X1 U22356 ( .A(n17039), .B(n2974), .Y(n16087) );
  OAI22XL U22357 ( .A0(n17060), .A1(n16087), .B0(n17061), .B1(n16008), .Y(
        n16092) );
  XNOR2X1 U22358 ( .A(n16289), .B(n3198), .Y(n16088) );
  OAI22X1 U22359 ( .A0(n16941), .A1(n16063), .B0(n16939), .B1(n16010), .Y(
        n16067) );
  XNOR2XL U22360 ( .A(n15968), .B(M3_mult_x_15_b_13_), .Y(n16089) );
  OAI22XL U22361 ( .A0(n16942), .A1(n16089), .B0(n16943), .B1(n16011), .Y(
        n16066) );
  OAI22X1 U22362 ( .A0(n16977), .A1(n16117), .B0(n3105), .B1(n16048), .Y(
        n16114) );
  XNOR2X1 U22363 ( .A(n3047), .B(n3196), .Y(n16116) );
  XNOR2XL U22364 ( .A(n16614), .B(n11495), .Y(n16107) );
  XNOR2X1 U22365 ( .A(n16614), .B(n3201), .Y(n16051) );
  OAI22XL U22366 ( .A0(n16942), .A1(n16020), .B0(n16943), .B1(n16126), .Y(
        n16146) );
  OAI22XL U22367 ( .A0(n17148), .A1(n12279), .B0(n3194), .B1(n11499), .Y(
        n16143) );
  CMPR32X1 U22368 ( .A(n11658), .B(n16022), .C(n16021), .CO(n16144), .S(n16023) );
  ADDFHX4 U22369 ( .A(n16025), .B(n16024), .CI(n16023), .CO(n16140), .S(n16018) );
  ADDFHX1 U22370 ( .A(n16028), .B(n16027), .CI(n16026), .CO(n16040), .S(n16035) );
  ADDFHX1 U22371 ( .A(n16031), .B(n16029), .CI(n16030), .CO(n16119), .S(n16039) );
  ADDFHX1 U22372 ( .A(n16056), .B(n16055), .CI(n16054), .CO(n16037), .S(n16073) );
  ADDFHX1 U22373 ( .A(n16062), .B(n16061), .CI(n16060), .CO(n16057), .S(n16787) );
  XNOR2X1 U22374 ( .A(n3203), .B(n16884), .Y(n16101) );
  OAI22XL U22375 ( .A0(n16941), .A1(n16101), .B0(n16939), .B1(n16063), .Y(
        n16112) );
  XNOR2X1 U22376 ( .A(n3022), .B(n3110), .Y(n16065) );
  OAI22XL U22377 ( .A0(n17092), .A1(n16065), .B0(n16317), .B1(n16064), .Y(
        n16111) );
  OAI22XL U22378 ( .A0(n17074), .A1(n16374), .B0(n16375), .B1(n16072), .Y(
        n16424) );
  ADDFHX4 U22379 ( .A(n16080), .B(n16079), .CI(n16078), .CO(n16852), .S(n16851) );
  ADDFHX1 U22380 ( .A(n16083), .B(n16082), .CI(n16081), .CO(n16076), .S(n16784) );
  XNOR2XL U22381 ( .A(n17039), .B(n11499), .Y(n16102) );
  OAI22XL U22382 ( .A0(n16942), .A1(n16115), .B0(n16943), .B1(n16089), .Y(
        n16104) );
  CMPR32X1 U22383 ( .A(n16094), .B(n16093), .C(n16092), .CO(n16097), .S(n16788) );
  OAI22XL U22384 ( .A0(n16941), .A1(n16373), .B0(n16939), .B1(n16101), .Y(
        n16443) );
  OAI22XL U22385 ( .A0(n16701), .A1(n16328), .B0(n16699), .B1(n16107), .Y(
        n16446) );
  XNOR2XL U22386 ( .A(n16289), .B(M3_mult_x_15_b_13_), .Y(n16331) );
  OAI22XL U22387 ( .A0(n16638), .A1(n16335), .B0(n16108), .B1(n16475), .Y(
        n16337) );
  OAI22XL U22388 ( .A0(n17074), .A1(n3212), .B0(n16375), .B1(n16109), .Y(
        n16336) );
  ADDFHX1 U22389 ( .A(n16112), .B(n16110), .CI(n16111), .CO(n16793), .S(n16814) );
  XNOR2X1 U22390 ( .A(n15968), .B(n3190), .Y(n16378) );
  OAI22XL U22391 ( .A0(n16942), .A1(n16378), .B0(n16688), .B1(n16115), .Y(
        n16431) );
  XNOR2X1 U22392 ( .A(n3199), .B(n3197), .Y(n16329) );
  OAI22XL U22393 ( .A0(n16977), .A1(n16329), .B0(n3105), .B1(n16117), .Y(
        n16429) );
  XNOR2XL U22394 ( .A(n3211), .B(M3_mult_x_15_b_13_), .Y(n16183) );
  XNOR2XL U22395 ( .A(n16289), .B(M3_mult_x_15_b_21_), .Y(n16165) );
  OAI22XL U22396 ( .A0(n17060), .A1(n16127), .B0(n17061), .B1(n16164), .Y(
        n16175) );
  XNOR2X1 U22397 ( .A(n17073), .B(M3_mult_x_15_b_9_), .Y(n16185) );
  OAI22XL U22398 ( .A0(n17074), .A1(n16128), .B0(n16375), .B1(n16185), .Y(
        n16174) );
  XNOR2X1 U22399 ( .A(n3199), .B(n3198), .Y(n16167) );
  XNOR2X1 U22400 ( .A(n3022), .B(n3197), .Y(n16184) );
  XNOR2X1 U22401 ( .A(n3203), .B(n3201), .Y(n16166) );
  CMPR32X1 U22402 ( .A(n12271), .B(n11658), .C(n16143), .CO(n16178), .S(n16145) );
  OAI22XL U22403 ( .A0(n17148), .A1(n11499), .B0(n17147), .B1(n3108), .Y(
        n16168) );
  CMPR32X1 U22404 ( .A(n16146), .B(n16145), .C(n16144), .CO(n16172), .S(n16141) );
  XNOR2X1 U22405 ( .A(n16289), .B(n3202), .Y(n16219) );
  OAI22XL U22406 ( .A0(n16867), .A1(n16166), .B0(n16939), .B1(n16200), .Y(
        n16222) );
  XNOR2XL U22407 ( .A(n3199), .B(n11495), .Y(n16202) );
  OAI22XL U22408 ( .A0(n16977), .A1(n16167), .B0(n3105), .B1(n16202), .Y(
        n16221) );
  CMPR32X1 U22409 ( .A(M3_mult_x_15_b_1_), .B(n12279), .C(n16168), .CO(n16220), 
        .S(n16177) );
  CMPR32X1 U22410 ( .A(n16176), .B(n16175), .C(n16174), .CO(n16199), .S(n16155) );
  OAI22XL U22411 ( .A0(n16701), .A1(n16614), .B0(n16699), .B1(n16605), .Y(
        n16205) );
  ADDFHX1 U22412 ( .A(n16182), .B(n16181), .CI(n16180), .CO(n16211), .S(n16158) );
  XNOR2X1 U22413 ( .A(n17073), .B(n16884), .Y(n16204) );
  OAI22XL U22414 ( .A0(n17074), .A1(n16185), .B0(n16375), .B1(n16204), .Y(
        n16216) );
  OAI22XL U22415 ( .A0(n16941), .A1(n16200), .B0(n16939), .B1(n16253), .Y(
        n16252) );
  XNOR2XL U22416 ( .A(n17039), .B(M3_mult_x_15_b_13_), .Y(n16241) );
  XNOR2X1 U22417 ( .A(n3199), .B(n3201), .Y(n16240) );
  OAI22XL U22418 ( .A0(n16893), .A1(n16202), .B0(n3105), .B1(n16240), .Y(
        n16250) );
  XNOR2X1 U22419 ( .A(n3022), .B(M3_mult_x_15_b_9_), .Y(n16242) );
  OAI22XL U22420 ( .A0(n17092), .A1(n16203), .B0(n16317), .B1(n16242), .Y(
        n16249) );
  XNOR2XL U22421 ( .A(n15968), .B(M3_mult_x_15_b_21_), .Y(n16238) );
  XNOR2X1 U22422 ( .A(n17073), .B(n3190), .Y(n16243) );
  OAI22XL U22423 ( .A0(n17074), .A1(n16204), .B0(n16375), .B1(n16243), .Y(
        n16247) );
  OAI22XL U22424 ( .A0(n17148), .A1(n3049), .B0(n17147), .B1(n3197), .Y(n16254) );
  ADDFHX1 U22425 ( .A(n16212), .B(n16211), .CI(n16210), .CO(n16260), .S(n16197) );
  ADDFHX1 U22426 ( .A(n16218), .B(n16217), .CI(n16216), .CO(n16234), .S(n16210) );
  XNOR2X1 U22427 ( .A(n3211), .B(n3198), .Y(n16239) );
  OAI2BB1XL U22428 ( .A0N(n16699), .A1N(n16701), .B0(n16614), .Y(n16235) );
  CMPR32X1 U22429 ( .A(n16237), .B(n16236), .C(n16235), .CO(n16292), .S(n16233) );
  OAI22XL U22430 ( .A0(n16942), .A1(n16238), .B0(n16943), .B1(n16288), .Y(
        n16272) );
  XNOR2XL U22431 ( .A(n3211), .B(n11495), .Y(n16287) );
  OAI22XL U22432 ( .A0(n16962), .A1(n16239), .B0(n16960), .B1(n16287), .Y(
        n16271) );
  XNOR2X1 U22433 ( .A(n3199), .B(n3196), .Y(n16280) );
  OAI22XL U22434 ( .A0(n16893), .A1(n16240), .B0(n3105), .B1(n16280), .Y(
        n16270) );
  XNOR2X1 U22435 ( .A(n17039), .B(n12701), .Y(n16275) );
  OAI22X1 U22436 ( .A0(n17060), .A1(n16241), .B0(n17061), .B1(n16275), .Y(
        n16286) );
  XNOR2X1 U22437 ( .A(n3022), .B(n16884), .Y(n16273) );
  OAI22X1 U22438 ( .A0(n17092), .A1(n16242), .B0(n16317), .B1(n16273), .Y(
        n16285) );
  XNOR2X1 U22439 ( .A(n5677), .B(n12561), .Y(n16274) );
  OAI22XL U22440 ( .A0(n17074), .A1(n16243), .B0(n16375), .B1(n16274), .Y(
        n16284) );
  CMPR32X1 U22441 ( .A(n16249), .B(n16248), .C(n16247), .CO(n16269), .S(n16256) );
  OAI22XL U22442 ( .A0(n16941), .A1(n16253), .B0(n16939), .B1(n16279), .Y(
        n16278) );
  CMPR32X1 U22443 ( .A(n11499), .B(n2974), .C(n16254), .CO(n16277), .S(n16231)
         );
  OAI22X1 U22444 ( .A0(n17148), .A1(n3197), .B0(n17147), .B1(
        M3_mult_x_15_n1682), .Y(n16282) );
  OAI22XL U22445 ( .A0(n3102), .A1(n16289), .B0(n16332), .B1(n16572), .Y(
        n16281) );
  CMPR32X1 U22446 ( .A(n16263), .B(n16262), .C(n16261), .CO(n16298), .S(n16295) );
  CMPR32X1 U22447 ( .A(n16269), .B(n16268), .C(n16267), .CO(n16304), .S(n16266) );
  CMPR32X1 U22448 ( .A(n16272), .B(n16271), .C(n16270), .CO(n16307), .S(n16291) );
  OAI22XL U22449 ( .A0(n17092), .A1(n16273), .B0(n16317), .B1(n16318), .Y(
        n16310) );
  XNOR2XL U22450 ( .A(n5677), .B(M3_mult_x_15_b_13_), .Y(n16320) );
  XNOR2X1 U22451 ( .A(n17039), .B(n3198), .Y(n16311) );
  OAI22XL U22452 ( .A0(n17060), .A1(n16275), .B0(n17061), .B1(n16311), .Y(
        n16308) );
  CMPR32X1 U22453 ( .A(n16278), .B(n16277), .C(n16276), .CO(n16305), .S(n16267) );
  XNOR2XL U22454 ( .A(n3203), .B(M3_mult_x_15_b_21_), .Y(n16312) );
  OAI22XL U22455 ( .A0(n16941), .A1(n16279), .B0(n16939), .B1(n16312), .Y(
        n16316) );
  OAI22XL U22456 ( .A0(n16893), .A1(n16280), .B0(n3105), .B1(n16313), .Y(
        n16315) );
  OAI22XL U22457 ( .A0(n17148), .A1(n5430), .B0(n17147), .B1(M3_mult_x_15_b_9_), .Y(n16321) );
  OAI22X1 U22458 ( .A0(n16942), .A1(n16288), .B0(n16943), .B1(n15968), .Y(
        n16323) );
  OAI2BB1XL U22459 ( .A0N(n16332), .A1N(n3102), .B0(n16289), .Y(n16322) );
  XNOR2X1 U22460 ( .A(n3203), .B(n3202), .Y(n16940) );
  XNOR2XL U22461 ( .A(n3199), .B(M3_mult_x_15_b_20_), .Y(n16976) );
  OAI22XL U22462 ( .A0(n16977), .A1(n16313), .B0(n3105), .B1(n16976), .Y(
        n16971) );
  XNOR2X1 U22463 ( .A(n3211), .B(n3196), .Y(n16961) );
  XNOR2X1 U22464 ( .A(n3022), .B(n12561), .Y(n16979) );
  OAI22XL U22465 ( .A0(n17092), .A1(n16318), .B0(n16317), .B1(n16979), .Y(
        n16957) );
  XNOR2X1 U22466 ( .A(n17073), .B(n12701), .Y(n16981) );
  CMPR32X1 U22467 ( .A(n3049), .B(n3197), .C(n16321), .CO(n16967), .S(n16314)
         );
  OAI22XL U22468 ( .A0(n16701), .A1(n16360), .B0(n16699), .B1(n16328), .Y(
        n16420) );
  XNOR2X1 U22469 ( .A(n3199), .B(M3_mult_x_15_b_6_), .Y(n16362) );
  XNOR2X1 U22470 ( .A(n16289), .B(n12561), .Y(n16333) );
  OAI22XL U22471 ( .A0(n3102), .A1(n16333), .B0(n16332), .B1(n16331), .Y(
        n16418) );
  OAI22XL U22472 ( .A0(n3102), .A1(n16351), .B0(n16332), .B1(n16333), .Y(
        n16392) );
  XNOR2X1 U22473 ( .A(M5_mult_x_15_n1), .B(n11495), .Y(n16341) );
  NOR2BX1 U22474 ( .AN(n3110), .B(n16375), .Y(n16340) );
  XNOR2X1 U22475 ( .A(n17039), .B(M3_mult_x_15_b_2_), .Y(n16377) );
  ADDHXL U22476 ( .A(n16337), .B(n16336), .CO(n16444), .S(n16423) );
  ADDFHX1 U22477 ( .A(n16340), .B(n16339), .CI(n16338), .CO(n16422), .S(n16390) );
  XNOR2X1 U22478 ( .A(n3203), .B(n3197), .Y(n16342) );
  XNOR2X1 U22479 ( .A(n3211), .B(n12279), .Y(n16347) );
  XNOR2XL U22480 ( .A(n3211), .B(n11499), .Y(n16383) );
  XNOR2X1 U22481 ( .A(n3047), .B(n3198), .Y(n16343) );
  XNOR2X1 U22482 ( .A(n3211), .B(M3_mult_x_15_b_1_), .Y(n16402) );
  OAI22XL U22483 ( .A0(n16962), .A1(n16402), .B0(n16960), .B1(n16348), .Y(
        n16398) );
  XNOR2X1 U22484 ( .A(n15968), .B(n3197), .Y(n16401) );
  XNOR2X1 U22485 ( .A(n15968), .B(M3_mult_x_15_n1682), .Y(n16353) );
  XNOR2X1 U22486 ( .A(n3047), .B(n12701), .Y(n16344) );
  XNOR2X1 U22487 ( .A(n3199), .B(n12279), .Y(n16404) );
  XNOR2XL U22488 ( .A(n3199), .B(n11499), .Y(n16350) );
  OAI22XL U22489 ( .A0(n16977), .A1(n16404), .B0(n3105), .B1(n16350), .Y(
        n16411) );
  OAI22X1 U22490 ( .A0(n16941), .A1(n16346), .B0(n16939), .B1(n16342), .Y(
        n16358) );
  OAI22XL U22491 ( .A0(n16701), .A1(n16345), .B0(n16699), .B1(n16361), .Y(
        n16356) );
  XNOR2X1 U22492 ( .A(n16614), .B(n3190), .Y(n16459) );
  XNOR2X1 U22493 ( .A(n3203), .B(n2974), .Y(n16409) );
  XNOR2X1 U22494 ( .A(n16289), .B(M3_mult_x_15_b_9_), .Y(n16410) );
  XNOR2X1 U22495 ( .A(n16289), .B(n16884), .Y(n16352) );
  OAI22XL U22496 ( .A0(n3102), .A1(n16410), .B0(n16332), .B1(n16352), .Y(
        n16412) );
  XNOR2X1 U22497 ( .A(n17039), .B(n3110), .Y(n16349) );
  XNOR2X1 U22498 ( .A(n3199), .B(n2974), .Y(n16363) );
  OAI22XL U22499 ( .A0(n16977), .A1(n16350), .B0(n3105), .B1(n16363), .Y(
        n16384) );
  XNOR2X1 U22500 ( .A(n4164), .B(M3_mult_x_15_b_9_), .Y(n16359) );
  ADDFHX1 U22501 ( .A(n16358), .B(n16357), .CI(n16356), .CO(n16369), .S(n16405) );
  XNOR2X1 U22502 ( .A(n15968), .B(n16884), .Y(n16379) );
  OAI22XL U22503 ( .A0(n16977), .A1(n16363), .B0(n3105), .B1(n16362), .Y(
        n16370) );
  ADDFHX1 U22504 ( .A(n16366), .B(n4764), .CI(n16364), .CO(n16421), .S(n16367)
         );
  ADDFHX1 U22505 ( .A(n16372), .B(n16371), .CI(n16370), .CO(n16437), .S(n16368) );
  OAI22XL U22506 ( .A0(n16962), .A1(n16383), .B0(n16960), .B1(n16382), .Y(
        n16438) );
  XNOR2X1 U22507 ( .A(M5_mult_x_15_n1), .B(n12701), .Y(n16462) );
  OAI22XL U22508 ( .A0(n16962), .A1(n16909), .B0(n16960), .B1(n16397), .Y(
        n16460) );
  XNOR2X1 U22509 ( .A(n15968), .B(M3_mult_x_15_b_6_), .Y(n16467) );
  XNOR2X1 U22510 ( .A(n3211), .B(n3110), .Y(n16403) );
  XNOR2X1 U22511 ( .A(n3199), .B(n12271), .Y(n16463) );
  OAI22XL U22512 ( .A0(n16977), .A1(n16463), .B0(n3105), .B1(n16404), .Y(
        n16470) );
  ADDFHX4 U22513 ( .A(n16407), .B(n16406), .CI(n16405), .CO(n16417), .S(n16479) );
  OAI22XL U22514 ( .A0(n16941), .A1(n16468), .B0(n16939), .B1(n16409), .Y(
        n16488) );
  OAI22XL U22515 ( .A0(n3102), .A1(n16474), .B0(n16332), .B1(n16410), .Y(
        n16487) );
  ADDFHX1 U22516 ( .A(n16423), .B(n16422), .CI(n16421), .CO(n16819), .S(n16447) );
  ADDFHX1 U22517 ( .A(n16426), .B(n16425), .CI(n16424), .CO(n16794), .S(n16799) );
  ADDFHX1 U22518 ( .A(n16431), .B(n16430), .CI(n16429), .CO(n16812), .S(n16797) );
  CMPR32X1 U22519 ( .A(n16446), .B(n16445), .C(n16444), .CO(n16815), .S(n16800) );
  CMPR22X1 U22520 ( .A(n16461), .B(n4805), .CO(n16466), .S(n16491) );
  XNOR2XL U22521 ( .A(M5_mult_x_15_n1), .B(M3_mult_x_15_b_13_), .Y(n16476) );
  OAI22X1 U22522 ( .A0(n16638), .A1(n16476), .B0(n16462), .B1(n16475), .Y(
        n16494) );
  XNOR2X1 U22523 ( .A(n3199), .B(M3_mult_x_15_b_1_), .Y(n16511) );
  OAI22XL U22524 ( .A0(n16977), .A1(n16511), .B0(n3105), .B1(n16463), .Y(
        n16493) );
  ADDFHX1 U22525 ( .A(n16466), .B(n16465), .CI(n16464), .CO(n16480), .S(n16503) );
  XNOR2X1 U22526 ( .A(n15968), .B(n2974), .Y(n16496) );
  OAI22XL U22527 ( .A0(n16942), .A1(n16496), .B0(n16688), .B1(n16467), .Y(
        n16501) );
  XNOR2X1 U22528 ( .A(n3203), .B(n12279), .Y(n16513) );
  XNOR2X1 U22529 ( .A(n3047), .B(n3190), .Y(n16497) );
  OAI22XL U22530 ( .A0(n16701), .A1(n16498), .B0(n16699), .B1(n16473), .Y(
        n16525) );
  XNOR2X1 U22531 ( .A(n16289), .B(n3197), .Y(n16510) );
  OAI22X1 U22532 ( .A0(n3102), .A1(n16510), .B0(n16332), .B1(n16474), .Y(
        n16524) );
  XNOR2X1 U22533 ( .A(M5_mult_x_15_n1), .B(n12561), .Y(n16518) );
  OAI22XL U22534 ( .A0(n16638), .A1(n16518), .B0(n16476), .B1(n16475), .Y(
        n16527) );
  OAI22XL U22535 ( .A0(n16893), .A1(n4796), .B0(n3105), .B1(n16477), .Y(n16526) );
  ADDFHX1 U22536 ( .A(n16486), .B(n16485), .CI(n16484), .CO(n16478), .S(n16563) );
  XNOR2X1 U22537 ( .A(n3047), .B(n16884), .Y(n16532) );
  OAI22XL U22538 ( .A0(n16701), .A1(n16533), .B0(n16699), .B1(n16498), .Y(
        n16514) );
  NAND2XL U22539 ( .A(n16777), .B(n16505), .Y(n16506) );
  OAI22XL U22540 ( .A0(n3102), .A1(n16531), .B0(n16332), .B1(n16510), .Y(
        n16522) );
  XNOR2X1 U22541 ( .A(n3199), .B(n3110), .Y(n16512) );
  OAI22XL U22542 ( .A0(n16977), .A1(n16512), .B0(n3105), .B1(n16511), .Y(
        n16521) );
  XNOR2X1 U22543 ( .A(n3203), .B(n12271), .Y(n16519) );
  OAI22XL U22544 ( .A0(n16941), .A1(n16519), .B0(n16939), .B1(n16513), .Y(
        n16520) );
  OAI22XL U22545 ( .A0(n16941), .A1(n16873), .B0(n16939), .B1(n16517), .Y(
        n16541) );
  XNOR2X1 U22546 ( .A(n3203), .B(M3_mult_x_15_b_1_), .Y(n16538) );
  OAI22XL U22547 ( .A0(n16941), .A1(n16538), .B0(n16939), .B1(n16519), .Y(
        n16528) );
  CMPR32X1 U22548 ( .A(n16522), .B(n16521), .C(n16520), .CO(n16554), .S(n16548) );
  ADDHXL U22549 ( .A(n16527), .B(n16526), .CO(n16523), .S(n16536) );
  ADDFHX1 U22550 ( .A(n16530), .B(n16529), .CI(n16528), .CO(n16535), .S(n16736) );
  XNOR2X1 U22551 ( .A(n16289), .B(n2974), .Y(n16537) );
  OAI22XL U22552 ( .A0(n3102), .A1(n16537), .B0(n16332), .B1(n16531), .Y(
        n16545) );
  XNOR2XL U22553 ( .A(n16289), .B(n11499), .Y(n16696) );
  OAI22XL U22554 ( .A0(n3102), .A1(n16696), .B0(n16332), .B1(n16537), .Y(
        n16707) );
  XNOR2X1 U22555 ( .A(n3203), .B(n3110), .Y(n16539) );
  XNOR2XL U22556 ( .A(n16614), .B(M3_mult_x_15_b_6_), .Y(n16698) );
  XNOR2XL U22557 ( .A(n15968), .B(M3_mult_x_15_b_2_), .Y(n16687) );
  ADDHXL U22558 ( .A(n16542), .B(n16541), .CO(n16737), .S(n16679) );
  CMPR32X1 U22559 ( .A(n16548), .B(n16547), .C(n16546), .CO(n16559), .S(n16733) );
  NAND2X1 U22560 ( .A(n16567), .B(n16770), .Y(n16772) );
  XNOR2X1 U22561 ( .A(n16289), .B(n12279), .Y(n16697) );
  OAI22XL U22562 ( .A0(n3102), .A1(n16577), .B0(n16332), .B1(n16697), .Y(
        n16692) );
  XNOR2X1 U22563 ( .A(n4164), .B(n3110), .Y(n16568) );
  XNOR2X1 U22564 ( .A(n15968), .B(M3_mult_x_15_b_1_), .Y(n16689) );
  XNOR2X1 U22565 ( .A(n16614), .B(n2974), .Y(n16700) );
  OAI22XL U22566 ( .A0(n16701), .A1(n16569), .B0(n16699), .B1(n16700), .Y(
        n16690) );
  XNOR2XL U22567 ( .A(n3047), .B(n2974), .Y(n16581) );
  OAI22XL U22568 ( .A0(n16701), .A1(n16584), .B0(n16699), .B1(n16569), .Y(
        n16586) );
  XNOR2X1 U22569 ( .A(M5_mult_x_15_n1), .B(M3_mult_x_15_b_6_), .Y(n16593) );
  XNOR2X1 U22570 ( .A(M5_mult_x_15_n1), .B(n3197), .Y(n16576) );
  OAI22XL U22571 ( .A0(n16638), .A1(n16593), .B0(n16576), .B1(n16475), .Y(
        n16592) );
  OAI22XL U22572 ( .A0(n3102), .A1(n16572), .B0(n16332), .B1(n16571), .Y(
        n16591) );
  XNOR2X1 U22573 ( .A(n3047), .B(n3197), .Y(n16703) );
  XNOR2X1 U22574 ( .A(M5_mult_x_15_n1), .B(M3_mult_x_15_b_9_), .Y(n16685) );
  XNOR2XL U22575 ( .A(n16289), .B(M3_mult_x_15_b_1_), .Y(n16582) );
  OAI22XL U22576 ( .A0(n3102), .A1(n16582), .B0(n16332), .B1(n16577), .Y(
        n16578) );
  XNOR2XL U22577 ( .A(n3047), .B(n11499), .Y(n16602) );
  XNOR2X1 U22578 ( .A(n16289), .B(n3110), .Y(n16583) );
  CMPR32X1 U22579 ( .A(n16587), .B(n16586), .C(n16585), .CO(n16721), .S(n16588) );
  NOR2XL U22580 ( .A(n16672), .B(n16671), .Y(n16675) );
  CMPR32X1 U22581 ( .A(n16590), .B(n16589), .C(n16588), .CO(n16671), .S(n16670) );
  ADDHXL U22582 ( .A(n16592), .B(n16591), .CO(n16585), .S(n16601) );
  XNOR2X1 U22583 ( .A(M5_mult_x_15_n1), .B(n2974), .Y(n16603) );
  NOR2XL U22584 ( .A(n16670), .B(n16669), .Y(n16598) );
  NOR2XL U22585 ( .A(n16675), .B(n16598), .Y(n16678) );
  XNOR2X1 U22586 ( .A(n3047), .B(n12279), .Y(n16613) );
  OAI22XL U22587 ( .A0(n16638), .A1(n16636), .B0(n16603), .B1(n16475), .Y(
        n16618) );
  NAND2BXL U22588 ( .AN(n3110), .B(n16614), .Y(n16604) );
  OAI22XL U22589 ( .A0(n16701), .A1(n16605), .B0(n16699), .B1(n16604), .Y(
        n16617) );
  NOR2XL U22590 ( .A(n16662), .B(n16661), .Y(n16609) );
  INVXL U22591 ( .A(n16609), .Y(n16665) );
  ADDHXL U22592 ( .A(n16618), .B(n16617), .CO(n16611), .S(n16648) );
  OR2X2 U22593 ( .A(n16660), .B(n16659), .Y(n16619) );
  NAND2XL U22594 ( .A(n16665), .B(n16619), .Y(n16668) );
  XNOR2X1 U22595 ( .A(M5_mult_x_15_n1), .B(n12271), .Y(n16628) );
  OAI22XL U22596 ( .A0(n16638), .A1(M3_mult_x_15_b_1_), .B0(n16628), .B1(
        n16475), .Y(n16624) );
  INVXL U22597 ( .A(n16624), .Y(n16627) );
  NAND2BX1 U22598 ( .AN(n2978), .B(M5_mult_x_15_n1), .Y(n16620) );
  INVXL U22599 ( .A(n16620), .Y(n16621) );
  NAND2XL U22600 ( .A(n16622), .B(n16621), .Y(n16626) );
  NAND2XL U22601 ( .A(n16624), .B(n16623), .Y(n16625) );
  OAI21XL U22602 ( .A0(n16627), .A1(n16626), .B0(n16625), .Y(n16635) );
  AOI21XL U22603 ( .A0(n16635), .A1(n16632), .B0(n6197), .Y(n16647) );
  OAI22XL U22604 ( .A0(n16638), .A1(n16637), .B0(n16636), .B1(n16475), .Y(
        n16652) );
  NOR2XL U22605 ( .A(n16644), .B(n16643), .Y(n16646) );
  NAND2XL U22606 ( .A(n16644), .B(n16643), .Y(n16645) );
  OAI21XL U22607 ( .A0(n16647), .A1(n16646), .B0(n16645), .Y(n16658) );
  CMPR32X1 U22608 ( .A(n16650), .B(n16649), .C(n16648), .CO(n16659), .S(n16656) );
  CMPR32X1 U22609 ( .A(n16653), .B(n16652), .C(n16651), .CO(n16655), .S(n16644) );
  AOI21XL U22610 ( .A0(n16658), .A1(n16654), .B0(n16657), .Y(n16667) );
  AND2X2 U22611 ( .A(n16662), .B(n16661), .Y(n16663) );
  AOI21XL U22612 ( .A0(n16665), .A1(n16664), .B0(n16663), .Y(n16666) );
  OAI21XL U22613 ( .A0(n16668), .A1(n16667), .B0(n16666), .Y(n16677) );
  NAND2XL U22614 ( .A(n16670), .B(n16669), .Y(n16674) );
  NAND2XL U22615 ( .A(n16672), .B(n16671), .Y(n16673) );
  OAI21XL U22616 ( .A0(n16675), .A1(n16674), .B0(n16673), .Y(n16676) );
  AOI21XL U22617 ( .A0(n16678), .A1(n16677), .B0(n16676), .Y(n16732) );
  CMPR32X1 U22618 ( .A(n16681), .B(n16680), .C(n16679), .CO(n16743), .S(n16750) );
  OAI22XL U22619 ( .A0(n16942), .A1(n16689), .B0(n16688), .B1(n16687), .Y(
        n16693) );
  OAI22XL U22620 ( .A0(n3102), .A1(n16697), .B0(n16332), .B1(n16696), .Y(
        n16710) );
  ADDFHX1 U22621 ( .A(n16719), .B(n16718), .CI(n16717), .CO(n16726), .S(n16725) );
  CMPR32X1 U22622 ( .A(n16722), .B(n16721), .C(n16720), .CO(n16724), .S(n16672) );
  OR2X2 U22623 ( .A(n16725), .B(n16724), .Y(n16723) );
  NAND2XL U22624 ( .A(n2998), .B(n16723), .Y(n16731) );
  AND2X2 U22625 ( .A(n16725), .B(n16724), .Y(n16729) );
  AND2X2 U22626 ( .A(n16727), .B(n16726), .Y(n16728) );
  AOI21X1 U22627 ( .A0(n2998), .A1(n16729), .B0(n16728), .Y(n16730) );
  CMPR32X1 U22628 ( .A(n16747), .B(n16746), .C(n16745), .CO(n16754), .S(n16753) );
  NOR2XL U22629 ( .A(n16753), .B(n16752), .Y(n16751) );
  NOR2XL U22630 ( .A(n16758), .B(n16751), .Y(n16760) );
  NAND2XL U22631 ( .A(n16753), .B(n16752), .Y(n16757) );
  NAND2XL U22632 ( .A(n16755), .B(n16754), .Y(n16756) );
  AND2X2 U22633 ( .A(n16768), .B(n16767), .Y(n16769) );
  ADDFHX4 U22634 ( .A(n16808), .B(n16807), .CI(n16806), .CO(n16848), .S(n16847) );
  XNOR2XL U22635 ( .A(n3199), .B(n3202), .Y(n16883) );
  OAI2BB1XL U22636 ( .A0N(n16939), .A1N(n16867), .B0(n3203), .Y(n16880) );
  XNOR2XL U22637 ( .A(n3211), .B(M3_mult_x_15_b_21_), .Y(n16869) );
  XNOR2X1 U22638 ( .A(n3022), .B(n12701), .Y(n16875) );
  OAI22XL U22639 ( .A0(n17092), .A1(n16875), .B0(n17099), .B1(n16871), .Y(
        n16878) );
  XNOR2XL U22640 ( .A(n5677), .B(n11495), .Y(n16874) );
  OAI22XL U22641 ( .A0(n17087), .A1(n16874), .B0(n16375), .B1(n16868), .Y(
        n16877) );
  XNOR2XL U22642 ( .A(n17039), .B(M3_mult_x_15_b_20_), .Y(n16888) );
  OAI22XL U22643 ( .A0(n17060), .A1(n16870), .B0(n17061), .B1(n16888), .Y(
        n16894) );
  OAI22XL U22644 ( .A0(n17148), .A1(n12561), .B0(n3194), .B1(
        M3_mult_x_15_b_13_), .Y(n16872) );
  OAI22XL U22645 ( .A0(n17148), .A1(M3_mult_x_15_b_13_), .B0(n3194), .B1(
        n12701), .Y(n16891) );
  OAI22XL U22646 ( .A0(n16977), .A1(n3199), .B0(n3105), .B1(n4796), .Y(n16890)
         );
  OAI22XL U22647 ( .A0(n16941), .A1(n3203), .B0(n16939), .B1(n16873), .Y(
        n16935) );
  XNOR2X1 U22648 ( .A(n17073), .B(n3198), .Y(n16980) );
  OAI22X1 U22649 ( .A0(n17074), .A1(n16980), .B0(n16375), .B1(n16874), .Y(
        n16946) );
  XNOR2XL U22650 ( .A(n3022), .B(M3_mult_x_15_b_13_), .Y(n16978) );
  XNOR2XL U22651 ( .A(n17039), .B(M3_mult_x_15_b_17_), .Y(n16937) );
  OAI22XL U22652 ( .A0(n17060), .A1(n16937), .B0(n17061), .B1(n16876), .Y(
        n16944) );
  CMPR32X1 U22653 ( .A(n16879), .B(n16878), .C(n16877), .CO(n16930), .S(n16949) );
  CMPR32X1 U22654 ( .A(n16882), .B(n16881), .C(n16880), .CO(n16931), .S(n16948) );
  XNOR2XL U22655 ( .A(n3199), .B(M3_mult_x_15_b_21_), .Y(n16975) );
  OAI22XL U22656 ( .A0(n16977), .A1(n16975), .B0(n3105), .B1(n16883), .Y(
        n16987) );
  OAI22XL U22657 ( .A0(n17148), .A1(n16884), .B0(n3194), .B1(n3190), .Y(n16963) );
  CMPR32X1 U22658 ( .A(n16887), .B(n16886), .C(n16885), .CO(n16902), .S(n16952) );
  XNOR2XL U22659 ( .A(n17039), .B(M3_mult_x_15_b_21_), .Y(n16904) );
  OAI22XL U22660 ( .A0(n17060), .A1(n16888), .B0(n17061), .B1(n16904), .Y(
        n16907) );
  CMPR32X1 U22661 ( .A(n12542), .B(n16891), .C(n16890), .CO(n16899), .S(n16885) );
  OAI2BB1XL U22662 ( .A0N(n3105), .A1N(n16893), .B0(n3199), .Y(n16910) );
  CMPR32X1 U22663 ( .A(n16902), .B(n16901), .C(n16900), .CO(n16914), .S(n16953) );
  XNOR2X1 U22664 ( .A(n17039), .B(n3202), .Y(n16923) );
  CMPR32X1 U22665 ( .A(n12561), .B(n12518), .C(n16908), .CO(n16918), .S(n16905) );
  CMPR32X1 U22666 ( .A(n16915), .B(n16914), .C(n16913), .CO(n17120), .S(n17117) );
  CMPR32X1 U22667 ( .A(n16918), .B(n16917), .C(n16916), .CO(n17034), .S(n16926) );
  ADDFHX1 U22668 ( .A(n16921), .B(n16920), .CI(n16919), .CO(n17049), .S(n16928) );
  CMPR32X1 U22669 ( .A(n3107), .B(n16925), .C(n16924), .CO(n17035), .S(n16917)
         );
  CMPR32X1 U22670 ( .A(n16928), .B(n16927), .C(n16926), .CO(n17032), .S(n16913) );
  CMPR32X1 U22671 ( .A(n16931), .B(n16930), .C(n16929), .CO(n16955), .S(n17010) );
  CMPR32X1 U22672 ( .A(n16934), .B(n16933), .C(n16932), .CO(n16951), .S(n17007) );
  OAI2BB1XL U22673 ( .A0N(n16943), .A1N(n16942), .B0(n4164), .Y(n16973) );
  CMPR32X1 U22674 ( .A(n16949), .B(n16948), .C(n16947), .CO(n16950), .S(n17005) );
  CMPR32X1 U22675 ( .A(n16952), .B(n16951), .C(n16950), .CO(n16954), .S(n17008) );
  OAI22XL U22676 ( .A0(n16962), .A1(n16961), .B0(n16960), .B1(n16959), .Y(
        n16990) );
  OAI22XL U22677 ( .A0(n17092), .A1(n16979), .B0(n17099), .B1(n16978), .Y(
        n16983) );
  OAI22XL U22678 ( .A0(n17074), .A1(n16981), .B0(n16319), .B1(n16980), .Y(
        n16982) );
  ADDFHX1 U22679 ( .A(n16983), .B(n16984), .CI(n16982), .CO(n17002), .S(n16994) );
  CMPR32X1 U22680 ( .A(n16987), .B(n16986), .C(n16985), .CO(n16947), .S(n17001) );
  ADDFHX1 U22681 ( .A(n16990), .B(n16989), .CI(n16988), .CO(n17000), .S(n16998) );
  CMPR32X1 U22682 ( .A(n17013), .B(n17012), .C(n17011), .CO(n17112), .S(n17110) );
  CMPR32X1 U22683 ( .A(n17031), .B(n17030), .C(n17029), .CO(n17111), .S(n17108) );
  CMPR32X1 U22684 ( .A(n17034), .B(n17033), .C(n17032), .CO(n17126), .S(n17119) );
  CMPR32X1 U22685 ( .A(n17037), .B(n17036), .C(n17035), .CO(n17052), .S(n17047) );
  OAI22X1 U22686 ( .A0(n17074), .A1(n17044), .B0(n16375), .B1(n17059), .Y(
        n17055) );
  OAI22XL U22687 ( .A0(n17092), .A1(n17045), .B0(n17099), .B1(n17058), .Y(
        n17054) );
  CMPR32X1 U22688 ( .A(n12701), .B(n3198), .C(n17046), .CO(n17053), .S(n17036)
         );
  CMPR32X1 U22689 ( .A(n17052), .B(n17051), .C(n17050), .CO(n17128), .S(n17125) );
  CMPR32X1 U22690 ( .A(n3043), .B(n17057), .C(n17056), .CO(n17076), .S(n17064)
         );
  XNOR2XL U22691 ( .A(n3022), .B(M3_mult_x_15_b_21_), .Y(n17071) );
  OAI22XL U22692 ( .A0(n17092), .A1(n17058), .B0(n17099), .B1(n17071), .Y(
        n17070) );
  CMPR32X1 U22693 ( .A(n17070), .B(n17069), .C(n17068), .CO(n17080), .S(n17075) );
  XNOR2X1 U22694 ( .A(n3022), .B(n3202), .Y(n17086) );
  CMPR32X1 U22695 ( .A(n3021), .B(n3201), .C(n17072), .CO(n17084), .S(n17077)
         );
  CMPR32X1 U22696 ( .A(n17077), .B(n17076), .C(n17075), .CO(n17078), .S(n17066) );
  CMPR32X1 U22697 ( .A(n5997), .B(n17082), .C(n17081), .CO(n17090), .S(n17083)
         );
  CMPR32X1 U22698 ( .A(n17085), .B(n17084), .C(n17083), .CO(n17089), .S(n17079) );
  CMPR32X1 U22699 ( .A(n17090), .B(n17089), .C(n17088), .CO(n17137), .S(n17134) );
  CMPR32X1 U22700 ( .A(n17095), .B(n17094), .C(n17093), .CO(n17096), .S(n17088) );
  CMPR32X1 U22701 ( .A(n17098), .B(n17097), .C(n17096), .CO(n17141), .S(n17136) );
  CMPR32X1 U22702 ( .A(n5960), .B(n17101), .C(n17100), .CO(n17102), .S(n17097)
         );
  NOR2X1 U22703 ( .A(n17141), .B(n17140), .Y(n17391) );
  CMPR32X1 U22704 ( .A(n17104), .B(n17103), .C(n17102), .CO(n17143), .S(n17140) );
  CMPR32X1 U22705 ( .A(M3_mult_x_15_b_20_), .B(M3_mult_x_15_b_21_), .C(n17105), 
        .CO(n17145), .S(n17103) );
  OR2X2 U22706 ( .A(n17143), .B(n17142), .Y(n17367) );
  OAI21XL U22707 ( .A0(n17348), .A1(n17342), .B0(n17349), .Y(n17121) );
  INVXL U22708 ( .A(n17310), .Y(n17354) );
  NAND2XL U22709 ( .A(n17130), .B(n17129), .Y(n17358) );
  INVXL U22710 ( .A(n17358), .Y(n17131) );
  AOI21XL U22711 ( .A0(n17354), .A1(n4634), .B0(n17131), .Y(n17132) );
  OAI21XL U22712 ( .A0(n17383), .A1(n17378), .B0(n17384), .Y(n17138) );
  CMPR32X1 U22713 ( .A(n5957), .B(n17146), .C(n17145), .CO(n17151), .S(n17142)
         );
  OAI21XL U22714 ( .A0(n26307), .A1(n15940), .B0(n17154), .Y(n17156) );
  OAI21XL U22715 ( .A0(n26292), .A1(n15940), .B0(n17157), .Y(n17159) );
  NOR2X1 U22716 ( .A(n17159), .B(n17158), .Y(n17397) );
  OAI21XL U22717 ( .A0(n26293), .A1(n17167), .B0(n17160), .Y(n17162) );
  OAI21XL U22718 ( .A0(n26300), .A1(n17167), .B0(n17166), .Y(n17169) );
  OAI21XL U22719 ( .A0(n26306), .A1(n17167), .B0(n17173), .Y(n17175) );
  CMPR32X1 U22720 ( .A(n18770), .B(n17186), .C(n17185), .CO(n17184), .S(n25132) );
  CMPR32X1 U22721 ( .A(n18773), .B(n17188), .C(n17187), .CO(n17195), .S(n25181) );
  CMPR32X1 U22722 ( .A(n18779), .B(n17192), .C(n17191), .CO(n17189), .S(n24360) );
  CMPR22X1 U22723 ( .A(n17397), .B(n18780), .CO(n17191), .S(n24359) );
  CMPR32X1 U22724 ( .A(n18783), .B(n17194), .C(n17193), .CO(n17185), .S(n25162) );
  CMPR32X1 U22725 ( .A(n18786), .B(n17196), .C(n17195), .CO(n17193), .S(n25107) );
  NAND4BXL U22726 ( .AN(n25132), .B(n17199), .C(n17198), .D(n17197), .Y(n17200) );
  NAND2XL U22727 ( .A(n17249), .B(n17254), .Y(n17219) );
  INVXL U22728 ( .A(n17253), .Y(n17217) );
  AOI21XL U22729 ( .A0(n17216), .A1(n17254), .B0(n17217), .Y(n17218) );
  INVXL U22730 ( .A(n17220), .Y(n17222) );
  NAND2XL U22731 ( .A(n17222), .B(n17221), .Y(n17223) );
  XNOR2X1 U22732 ( .A(n17224), .B(n17223), .Y(n17452) );
  INVX1 U22733 ( .A(n17241), .Y(n17304) );
  INVXL U22734 ( .A(n17231), .Y(n17233) );
  NAND2XL U22735 ( .A(n17238), .B(n17303), .Y(n17244) );
  OAI21XL U22736 ( .A0(n3158), .A1(n17237), .B0(n17307), .Y(n17240) );
  INVXL U22737 ( .A(n17245), .Y(n17247) );
  INVXL U22738 ( .A(n17249), .Y(n17251) );
  NAND2XL U22739 ( .A(n17254), .B(n17253), .Y(n17255) );
  XNOR2X1 U22740 ( .A(n17256), .B(n17255), .Y(n17450) );
  INVXL U22741 ( .A(n17258), .Y(n17259) );
  INVXL U22742 ( .A(n17260), .Y(n17262) );
  NAND2XL U22743 ( .A(n17262), .B(n17261), .Y(n17263) );
  OAI21XL U22744 ( .A0(n17284), .A1(n18818), .B0(n17286), .Y(n17267) );
  OAI21XL U22745 ( .A0(M3_U4_U1_enc_tree_2__4__16_), .A1(
        M5_U3_U1_enc_tree_2__4__16_), .B0(n17267), .Y(n17271) );
  NAND2XL U22746 ( .A(n17303), .B(n17297), .Y(n17298) );
  INVXL U22747 ( .A(n17295), .Y(n17296) );
  INVXL U22748 ( .A(n17299), .Y(n17301) );
  NAND2XL U22749 ( .A(n17303), .B(n17236), .Y(n17306) );
  NAND2X1 U22750 ( .A(n3161), .B(n17307), .Y(n17308) );
  INVX1 U22751 ( .A(n17309), .Y(n17352) );
  INVXL U22752 ( .A(n17311), .Y(n17319) );
  NAND2XL U22753 ( .A(n17335), .B(n17339), .Y(n17323) );
  NOR2XL U22754 ( .A(n17319), .B(n17323), .Y(n17341) );
  INVXL U22755 ( .A(n17320), .Y(n17334) );
  AOI21XL U22756 ( .A0(n17334), .A1(n17339), .B0(n17321), .Y(n17322) );
  OAI21XL U22757 ( .A0(n17324), .A1(n17323), .B0(n17322), .Y(n17345) );
  INVXL U22758 ( .A(n17345), .Y(n17325) );
  NAND2XL U22759 ( .A(n17311), .B(n17328), .Y(n17330) );
  NAND2XL U22760 ( .A(n17311), .B(n17335), .Y(n17337) );
  AOI21XL U22761 ( .A0(n17312), .A1(n17335), .B0(n17334), .Y(n17336) );
  INVXL U22762 ( .A(n17342), .Y(n17343) );
  AOI21XL U22763 ( .A0(n17345), .A1(n17344), .B0(n17343), .Y(n17346) );
  INVXL U22764 ( .A(n17348), .Y(n17350) );
  NAND2XL U22765 ( .A(n17353), .B(n17355), .Y(n17357) );
  INVXL U22766 ( .A(n17360), .Y(n17361) );
  NAND2XL U22767 ( .A(n3149), .B(n17363), .Y(n17365) );
  INVXL U22768 ( .A(n17370), .Y(n17374) );
  INVX1 U22769 ( .A(n17376), .Y(n17380) );
  NAND2XL U22770 ( .A(n17377), .B(n17380), .Y(n17382) );
  INVXL U22771 ( .A(n17388), .Y(n17389) );
  NOR2XL U22772 ( .A(n17434), .B(n4855), .Y(n17424) );
  XOR2X1 U22773 ( .A(n17426), .B(n17425), .Y(n17439) );
  NAND2XL U22774 ( .A(n3357), .B(n17428), .Y(n17429) );
  INVXL U22775 ( .A(n17441), .Y(n17442) );
  NAND2XL U22776 ( .A(n20735), .B(n17442), .Y(n20333) );
  NAND2X1 U22777 ( .A(n17448), .B(n5336), .Y(n17449) );
  NOR2XL U22778 ( .A(n20340), .B(n20341), .Y(n17451) );
  INVXL U22779 ( .A(n17452), .Y(n17453) );
  XOR2X1 U22780 ( .A(n17454), .B(n17453), .Y(n20343) );
  OAI21XL U22781 ( .A0(n3045), .A1(n25912), .B0(n17460), .Y(n17461) );
  INVXL U22782 ( .A(n17469), .Y(n17472) );
  INVXL U22783 ( .A(n17470), .Y(n17471) );
  AOI22X1 U22784 ( .A0(n5480), .A1(sigma11[19]), .B0(in_valid_t), .B1(w2[51]), 
        .Y(n17476) );
  OAI21X2 U22785 ( .A0(n25813), .A1(n26254), .B0(n17476), .Y(M4_a_19_) );
  NAND2X1 U22786 ( .A(n3132), .B(n17487), .Y(n17488) );
  NAND2X1 U22787 ( .A(n3132), .B(n17489), .Y(n17490) );
  CLKINVX3 U22788 ( .A(n20993), .Y(n23534) );
  NAND2X2 U22789 ( .A(n17501), .B(n17491), .Y(n18483) );
  BUFX8 U22790 ( .A(n18483), .Y(n18522) );
  CLKINVX8 U22791 ( .A(n18467), .Y(n18468) );
  XNOR2X1 U22792 ( .A(n18468), .B(n3190), .Y(n17509) );
  BUFX8 U22793 ( .A(n17937), .Y(n18242) );
  XNOR2X1 U22794 ( .A(n3206), .B(n3202), .Y(n17519) );
  XOR2X1 U22795 ( .A(M4_a_4_), .B(M4_a_5_), .Y(n17492) );
  NAND2X2 U22796 ( .A(n17492), .B(n18141), .Y(n17861) );
  INVX2 U22797 ( .A(M4_a_5_), .Y(n18142) );
  XNOR2XL U22798 ( .A(n18150), .B(M3_mult_x_15_b_21_), .Y(n17503) );
  XNOR2X1 U22799 ( .A(n18118), .B(M5_b_18_), .Y(n17517) );
  XNOR2X1 U22800 ( .A(n18118), .B(n3048), .Y(n17505) );
  INVX4 U22801 ( .A(M4_a_17_), .Y(n18603) );
  CLKBUFX8 U22802 ( .A(n17493), .Y(n18625) );
  XNOR2X1 U22803 ( .A(n18604), .B(M3_mult_x_15_b_9_), .Y(n17507) );
  XNOR2X1 U22804 ( .A(n18638), .B(n3049), .Y(n17528) );
  BUFX4 U22805 ( .A(n18653), .Y(n17872) );
  XNOR2X1 U22806 ( .A(n18638), .B(n3197), .Y(n17496) );
  OAI22X1 U22807 ( .A0(n18652), .A1(n17528), .B0(n17872), .B1(n17496), .Y(
        n17530) );
  XNOR2X1 U22808 ( .A(n18453), .B(n18611), .Y(n17510) );
  XNOR2X1 U22809 ( .A(n25883), .B(n2974), .Y(n17553) );
  XNOR2X1 U22810 ( .A(n25883), .B(n3049), .Y(n17511) );
  OAI22XL U22811 ( .A0(n18652), .A1(n17496), .B0(n17872), .B1(n17500), .Y(
        n17497) );
  ADDFHX1 U22812 ( .A(n17499), .B(n17498), .CI(n17497), .CO(n17612), .S(n17575) );
  XNOR2X1 U22813 ( .A(n18638), .B(M3_mult_x_15_b_9_), .Y(n17638) );
  OAI22X1 U22814 ( .A0(n18652), .A1(n17500), .B0(n17872), .B1(n17638), .Y(
        n17632) );
  INVX2 U22815 ( .A(M4_a_9_), .Y(n18110) );
  INVX8 U22816 ( .A(n18110), .Y(n18503) );
  XNOR2X1 U22817 ( .A(n18503), .B(n3048), .Y(n17621) );
  XNOR2X1 U22818 ( .A(n18150), .B(n3202), .Y(n17502) );
  OAI22X1 U22819 ( .A0(n17861), .A1(n17502), .B0(n18141), .B1(n18150), .Y(
        n17617) );
  OAI22XL U22820 ( .A0(n18107), .A1(n17504), .B0(n17902), .B1(n17620), .Y(
        n17616) );
  XNOR2X1 U22821 ( .A(n18500), .B(n3198), .Y(n17516) );
  BUFX4 U22822 ( .A(n18501), .Y(n18429) );
  OAI22XL U22823 ( .A0(n18083), .A1(n17516), .B0(n18429), .B1(n17558), .Y(
        n17568) );
  OAI22XL U22824 ( .A0(n18239), .A1(n17503), .B0(n18141), .B1(n17502), .Y(
        n17567) );
  XNOR2X1 U22825 ( .A(n18453), .B(n3198), .Y(n17623) );
  OAI22X1 U22826 ( .A0(n18659), .A1(n17511), .B0(n17832), .B1(n17637), .Y(
        n17640) );
  OAI2BB1XL U22827 ( .A0N(n18168), .A1N(n17937), .B0(n3206), .Y(n17639) );
  XNOR2X1 U22828 ( .A(n18503), .B(n3021), .Y(n17513) );
  OAI22XL U22829 ( .A0(n18111), .A1(n17538), .B0(n18504), .B1(n17513), .Y(
        n17585) );
  BUFX3 U22830 ( .A(n17962), .Y(n18223) );
  XNOR2X1 U22831 ( .A(n18503), .B(n3201), .Y(n17521) );
  OAI22XL U22832 ( .A0(n18111), .A1(n17513), .B0(n18504), .B1(n17521), .Y(
        n17526) );
  ADDFHX1 U22833 ( .A(n2978), .B(n17515), .CI(n17514), .CO(n17525), .S(n17583)
         );
  XNOR2X1 U22834 ( .A(n25883), .B(M3_mult_x_15_b_2_), .Y(n17586) );
  XNOR2X1 U22835 ( .A(n25883), .B(M3_mult_x_15_b_3_), .Y(n17527) );
  OAI22X1 U22836 ( .A0(n18659), .A1(n17586), .B0(n17832), .B1(n17527), .Y(
        n17588) );
  XNOR2X1 U22837 ( .A(n18638), .B(n2974), .Y(n17529) );
  XNOR2X1 U22838 ( .A(n3206), .B(M3_mult_x_15_b_21_), .Y(n17536) );
  OAI22X1 U22839 ( .A0(n18242), .A1(n17536), .B0(n18168), .B1(n17519), .Y(
        n17548) );
  XNOR2X1 U22840 ( .A(n18150), .B(n3048), .Y(n17537) );
  OAI22XL U22841 ( .A0(n18239), .A1(n17537), .B0(n18141), .B1(n17520), .Y(
        n17547) );
  ADDFHX1 U22842 ( .A(n11658), .B(n17523), .CI(n17522), .CO(n17560), .S(n17524) );
  ADDFHX1 U22843 ( .A(n17526), .B(n17525), .CI(n17524), .CO(n17556), .S(n17593) );
  XNOR2X1 U22844 ( .A(n18453), .B(n3190), .Y(n17535) );
  XNOR2XL U22845 ( .A(n25883), .B(n11499), .Y(n17554) );
  OAI22XL U22846 ( .A0(n18652), .A1(n17529), .B0(n17872), .B1(n17528), .Y(
        n17542) );
  XNOR2XL U22847 ( .A(n18453), .B(M4_mult_x_15_n1680), .Y(n17654) );
  XNOR2X1 U22848 ( .A(n18150), .B(n3196), .Y(n17657) );
  OAI22XL U22849 ( .A0(n18239), .A1(n17657), .B0(n18141), .B1(n17537), .Y(
        n17662) );
  ADDFHX1 U22850 ( .A(n17544), .B(n17543), .CI(n17542), .CO(n17546), .S(n17597) );
  ADDFHX1 U22851 ( .A(n17549), .B(n17548), .CI(n17547), .CO(n17571), .S(n17595) );
  OAI22X1 U22852 ( .A0(n18659), .A1(n17554), .B0(n17832), .B1(n17553), .Y(
        n17563) );
  XNOR2X1 U22853 ( .A(n18500), .B(n3201), .Y(n17622) );
  OAI22XL U22854 ( .A0(n18083), .A1(n17558), .B0(n18429), .B1(n17622), .Y(
        n17635) );
  OAI22XL U22855 ( .A0(n18721), .A1(n11499), .B0(n17512), .B1(n3108), .Y(
        n17624) );
  ADDFHX1 U22856 ( .A(n17562), .B(n17561), .CI(n17560), .CO(n17629), .S(n17557) );
  ADDFHX1 U22857 ( .A(n17564), .B(n17563), .CI(M4_U3_U1_or2_inv_0__30_), .CO(
        n17574), .S(n17569) );
  ADDFHX1 U22858 ( .A(n17571), .B(n17570), .CI(n17569), .CO(n17580), .S(n17651) );
  ADDFHX1 U22859 ( .A(n17574), .B(n17573), .CI(n17572), .CO(n17628), .S(n17579) );
  ADDFHX1 U22860 ( .A(n17577), .B(n17576), .CI(n17575), .CO(n17644), .S(n17578) );
  ADDFHX1 U22861 ( .A(n17580), .B(n17579), .CI(n17578), .CO(n17625), .S(n17650) );
  XNOR2X1 U22862 ( .A(n18604), .B(n3049), .Y(n17601) );
  XNOR2X1 U22863 ( .A(n18468), .B(n5430), .Y(n17600) );
  OAI22XL U22864 ( .A0(n18522), .A1(n17600), .B0(n3195), .B1(n17582), .Y(
        n17659) );
  ADDFHX1 U22865 ( .A(n17589), .B(n17588), .CI(n17587), .CO(n17596), .S(n17669) );
  XNOR2X1 U22866 ( .A(n18468), .B(n3197), .Y(n17678) );
  XNOR2X1 U22867 ( .A(n18638), .B(M3_mult_x_15_b_3_), .Y(n17674) );
  OAI22XL U22868 ( .A0(n18624), .A1(n17693), .B0(n18625), .B1(n17601), .Y(
        n17699) );
  XNOR2XL U22869 ( .A(n18503), .B(M3_mult_x_15_b_13_), .Y(n17695) );
  XNOR2X1 U22870 ( .A(n18500), .B(M3_mult_x_15_b_11_), .Y(n17671) );
  XNOR2X1 U22871 ( .A(n18118), .B(n3198), .Y(n17694) );
  OAI22XL U22872 ( .A0(n18107), .A1(n17694), .B0(n17902), .B1(n17603), .Y(
        n17675) );
  NAND2BX1 U22873 ( .AN(n2978), .B(n25883), .Y(n17606) );
  XNOR2X1 U22874 ( .A(n3196), .B(n3206), .Y(n17718) );
  XNOR2X1 U22875 ( .A(n18150), .B(n3201), .Y(n17658) );
  NOR2X1 U22876 ( .A(n18406), .B(n18405), .Y(n18907) );
  OAI22XL U22877 ( .A0(n18083), .A1(n17622), .B0(n18429), .B1(n17746), .Y(
        n17738) );
  XNOR2X1 U22878 ( .A(n18453), .B(n3021), .Y(n17750) );
  CMPR32X1 U22879 ( .A(n17635), .B(n17634), .C(n17633), .CO(n17799), .S(n17630) );
  XNOR2X1 U22880 ( .A(n18468), .B(n18611), .Y(n17734) );
  XNOR2XL U22881 ( .A(n18638), .B(M4_mult_x_15_n1680), .Y(n17745) );
  OAI22X1 U22882 ( .A0(n18721), .A1(n3108), .B0(n17512), .B1(n3049), .Y(n17728) );
  OAI22XL U22883 ( .A0(n18239), .A1(n18150), .B0(n18141), .B1(n18142), .Y(
        n17727) );
  ADDFHX1 U22884 ( .A(n17641), .B(n17640), .CI(n17639), .CO(n17764), .S(n17613) );
  ADDFHX1 U22885 ( .A(n17650), .B(n17649), .CI(n17648), .CO(n18405), .S(n18403) );
  OAI22XL U22886 ( .A0(n18541), .A1(n17655), .B0(n5893), .B1(n17654), .Y(
        n17698) );
  OAI22XL U22887 ( .A0(n17861), .A1(n17658), .B0(n18141), .B1(n17657), .Y(
        n17696) );
  ADDFHX1 U22888 ( .A(n17664), .B(n17663), .CI(n17662), .CO(n17599), .S(n17682) );
  XNOR2XL U22889 ( .A(n25883), .B(n2978), .Y(n17673) );
  OAI22X1 U22890 ( .A0(n18659), .A1(n17673), .B0(n17832), .B1(n17672), .Y(
        n17722) );
  OAI22XL U22891 ( .A0(n18652), .A1(n17681), .B0(n17872), .B1(n17674), .Y(
        n17721) );
  CMPR32X1 U22892 ( .A(n17677), .B(n17676), .C(n17675), .CO(n17703), .S(n18342) );
  XNOR2X1 U22893 ( .A(n18468), .B(n3049), .Y(n17709) );
  OAI22XL U22894 ( .A0(n18522), .A1(n17709), .B0(n3195), .B1(n17678), .Y(
        n18346) );
  NOR2BX1 U22895 ( .AN(n2978), .B(n17832), .Y(n17869) );
  XNOR2X1 U22896 ( .A(n18006), .B(n3048), .Y(n17715) );
  XNOR2XL U22897 ( .A(n18604), .B(n11499), .Y(n17708) );
  XNOR2X1 U22898 ( .A(n18118), .B(n18611), .Y(n17714) );
  OAI22X1 U22899 ( .A0(n18107), .A1(n17714), .B0(n17902), .B1(n17694), .Y(
        n17711) );
  XNOR2X1 U22900 ( .A(n18503), .B(n12561), .Y(n17717) );
  OAI22XL U22901 ( .A0(n18111), .A1(n17717), .B0(n18504), .B1(n17695), .Y(
        n17710) );
  XNOR2X1 U22902 ( .A(n18604), .B(M3_mult_x_15_b_3_), .Y(n17874) );
  XNOR2X1 U22903 ( .A(n18468), .B(n2974), .Y(n17896) );
  OAI22XL U22904 ( .A0(n18522), .A1(n17896), .B0(n3195), .B1(n17709), .Y(
        n17926) );
  XNOR2X1 U22905 ( .A(n18150), .B(n3198), .Y(n17860) );
  OAI22XL U22906 ( .A0(n18239), .A1(n17860), .B0(n18141), .B1(n17713), .Y(
        n17931) );
  XNOR2XL U22907 ( .A(n18118), .B(M3_mult_x_15_b_13_), .Y(n17863) );
  OAI22XL U22908 ( .A0(n18107), .A1(n17863), .B0(n17902), .B1(n17714), .Y(
        n17930) );
  XNOR2X1 U22909 ( .A(n18006), .B(n3196), .Y(n17866) );
  NAND2BX1 U22910 ( .AN(n2978), .B(n18638), .Y(n17716) );
  OAI22XL U22911 ( .A0(n18652), .A1(n18637), .B0(n17872), .B1(n17716), .Y(
        n17864) );
  XNOR2X1 U22912 ( .A(n18503), .B(n3190), .Y(n17892) );
  XNOR2X1 U22913 ( .A(n3206), .B(n3201), .Y(n17894) );
  OAI22X1 U22914 ( .A0(n17937), .A1(n17894), .B0(n18168), .B1(n17718), .Y(
        n17877) );
  XNOR2X1 U22915 ( .A(n18453), .B(n3197), .Y(n17862) );
  OAI22XL U22916 ( .A0(n18721), .A1(n3049), .B0(n17512), .B1(n3197), .Y(n17752) );
  ADDFHX1 U22917 ( .A(n17733), .B(n17732), .CI(n17731), .CO(n17771), .S(n17762) );
  OAI2BB1XL U22918 ( .A0N(n18141), .A1N(n17861), .B0(n18150), .Y(n17739) );
  CMPR32X1 U22919 ( .A(n17738), .B(n17737), .C(n17736), .CO(n17770), .S(n17767) );
  XNOR2X1 U22920 ( .A(n18503), .B(n3202), .Y(n17791) );
  XNOR2X1 U22921 ( .A(n18468), .B(n3021), .Y(n17790) );
  XNOR2X1 U22922 ( .A(n18453), .B(n3201), .Y(n17749) );
  XNOR2X1 U22923 ( .A(n18453), .B(n3196), .Y(n17784) );
  XNOR2XL U22924 ( .A(n18604), .B(M3_mult_x_15_b_13_), .Y(n17747) );
  XNOR2X1 U22925 ( .A(n25883), .B(M3_mult_x_15_b_9_), .Y(n17742) );
  XNOR2XL U22926 ( .A(n18638), .B(M3_mult_x_15_b_11_), .Y(n17744) );
  XNOR2XL U22927 ( .A(n18638), .B(M3_mult_x_15_b_12_), .Y(n17778) );
  OAI22XL U22928 ( .A0(n18652), .A1(n17744), .B0(n17872), .B1(n17778), .Y(
        n17787) );
  OAI22XL U22929 ( .A0(n18652), .A1(n17745), .B0(n17872), .B1(n17744), .Y(
        n17756) );
  XNOR2X1 U22930 ( .A(n18500), .B(n3048), .Y(n17751) );
  OAI22XL U22931 ( .A0(n18083), .A1(n17746), .B0(n18429), .B1(n17751), .Y(
        n17755) );
  OAI22XL U22932 ( .A0(n18624), .A1(n17748), .B0(n18625), .B1(n17747), .Y(
        n17754) );
  OAI22XL U22933 ( .A0(n18541), .A1(n17750), .B0(n18539), .B1(n17749), .Y(
        n17753) );
  OAI22XL U22934 ( .A0(n18083), .A1(n17751), .B0(n18429), .B1(n17783), .Y(
        n17782) );
  CMPR32X1 U22935 ( .A(n11499), .B(n2974), .C(n17752), .CO(n17781), .S(n17761)
         );
  OAI22XL U22936 ( .A0(n18107), .A1(n18118), .B0(n17902), .B1(n18106), .Y(
        n17785) );
  CMPR32X1 U22937 ( .A(n17758), .B(n17757), .C(n17756), .CO(n17774), .S(n17802) );
  NAND2XL U22938 ( .A(n17764), .B(n17763), .Y(n17765) );
  OAI22XL U22939 ( .A0(n18652), .A1(n17778), .B0(n17872), .B1(n17834), .Y(
        n17823) );
  XNOR2X1 U22940 ( .A(n18604), .B(n3198), .Y(n17825) );
  OAI22XL U22941 ( .A0(n18624), .A1(n17779), .B0(n18625), .B1(n17825), .Y(
        n17822) );
  OAI22XL U22942 ( .A0(n18083), .A1(n17783), .B0(n18429), .B1(n17826), .Y(
        n17830) );
  XNOR2X1 U22943 ( .A(n18453), .B(n3048), .Y(n17827) );
  OAI22XL U22944 ( .A0(n18541), .A1(n17784), .B0(n18539), .B1(n17827), .Y(
        n17829) );
  OAI22XL U22945 ( .A0(n18721), .A1(n5430), .B0(n17512), .B1(M3_mult_x_15_b_9_), .Y(n17835) );
  ADDFHX1 U22946 ( .A(n16283), .B(n17786), .CI(n17785), .CO(n17841), .S(n17780) );
  XNOR2X1 U22947 ( .A(n18468), .B(n3201), .Y(n17831) );
  OAI22XL U22948 ( .A0(n18483), .A1(n17790), .B0(n3195), .B1(n17831), .Y(
        n17838) );
  OAI2BB1XL U22949 ( .A0N(n17902), .A1N(n18107), .B0(n18118), .Y(n17836) );
  ADDFHX1 U22950 ( .A(n17794), .B(n17793), .CI(n17792), .CO(n17813), .S(n17795) );
  CMPR32X1 U22951 ( .A(n17803), .B(n17802), .C(n17801), .CO(n17808), .S(n17846) );
  ADDFHX1 U22952 ( .A(n17809), .B(n17808), .CI(n17807), .CO(n17811), .S(n17857) );
  XNOR2X1 U22953 ( .A(n18500), .B(n3202), .Y(n18502) );
  OAI22X1 U22954 ( .A0(n18083), .A1(n17826), .B0(n18429), .B1(n18502), .Y(
        n18533) );
  OAI22XL U22955 ( .A0(n18541), .A1(n17827), .B0(n18539), .B1(n18540), .Y(
        n18532) );
  CMPR32X1 U22956 ( .A(n17830), .B(n17829), .C(n17828), .CO(n18554), .S(n17815) );
  XNOR2X1 U22957 ( .A(n18468), .B(n3196), .Y(n18521) );
  OAI22XL U22958 ( .A0(n18522), .A1(n17831), .B0(n3195), .B1(n18521), .Y(
        n18519) );
  XNOR2X1 U22959 ( .A(n25883), .B(n12561), .Y(n18543) );
  CMPR32X1 U22960 ( .A(n3049), .B(n3197), .C(n17835), .CO(n18528), .S(n17828)
         );
  OAI22XL U22961 ( .A0(n18111), .A1(n18503), .B0(n18504), .B1(n18110), .Y(
        n18524) );
  ADDFHX1 U22962 ( .A(n17850), .B(n17849), .CI(n17848), .CO(n17854), .S(n17851) );
  XNOR2X1 U22963 ( .A(n18150), .B(n18611), .Y(n17881) );
  OAI22XL U22964 ( .A0(n17861), .A1(n17881), .B0(n18141), .B1(n17860), .Y(
        n17917) );
  XNOR2X1 U22965 ( .A(n18453), .B(n3049), .Y(n17882) );
  OAI22XL U22966 ( .A0(n18107), .A1(n17906), .B0(n17902), .B1(n17863), .Y(
        n17915) );
  ADDHXL U22967 ( .A(n17865), .B(n17864), .CO(n17929), .S(n17922) );
  NOR2BX1 U22968 ( .AN(n2978), .B(n17872), .Y(n17911) );
  XNOR2X1 U22969 ( .A(n18604), .B(M3_mult_x_15_b_2_), .Y(n17875) );
  OAI22XL U22970 ( .A0(n18624), .A1(n17899), .B0(n18625), .B1(n17875), .Y(
        n17909) );
  XNOR2X1 U22971 ( .A(n18468), .B(M3_mult_x_15_b_3_), .Y(n17898) );
  XNOR2XL U22972 ( .A(n18468), .B(n11499), .Y(n17897) );
  OAI22X1 U22973 ( .A0(n18522), .A1(n17898), .B0(n3195), .B1(n17897), .Y(
        n17884) );
  XNOR2X1 U22974 ( .A(n3206), .B(n3198), .Y(n17880) );
  XNOR2X1 U22975 ( .A(n3206), .B(n3021), .Y(n17895) );
  OAI22XL U22976 ( .A0(n18242), .A1(n17880), .B0(n18168), .B1(n17895), .Y(
        n17883) );
  ADDFHX1 U22977 ( .A(n17869), .B(n17868), .CI(n17867), .CO(n18344), .S(n18349) );
  OAI22XL U22978 ( .A0(n18624), .A1(n17875), .B0(n18625), .B1(n17874), .Y(
        n17889) );
  XNOR2X1 U22979 ( .A(n3206), .B(n18611), .Y(n17936) );
  OAI22X1 U22980 ( .A0(n18242), .A1(n17936), .B0(n18168), .B1(n17880), .Y(
        n17940) );
  XNOR2XL U22981 ( .A(n18503), .B(M3_mult_x_15_b_9_), .Y(n17903) );
  XNOR2X1 U22982 ( .A(n18453), .B(n2974), .Y(n17901) );
  ADDFHX1 U22983 ( .A(n17885), .B(n17884), .CI(n17883), .CO(n17920), .S(n17950) );
  ADDFHX1 U22984 ( .A(n17886), .B(n17887), .CI(n17888), .CO(n17914), .S(n17951) );
  OAI22XL U22985 ( .A0(n18111), .A1(n17893), .B0(n18504), .B1(n17892), .Y(
        n17925) );
  OAI22X1 U22986 ( .A0(n18242), .A1(n17895), .B0(n18168), .B1(n17894), .Y(
        n17924) );
  OAI22XL U22987 ( .A0(n18522), .A1(n17897), .B0(n3195), .B1(n17896), .Y(
        n17923) );
  OAI22XL U22988 ( .A0(n18522), .A1(n17935), .B0(n3195), .B1(n17898), .Y(
        n17946) );
  XNOR2XL U22989 ( .A(n18453), .B(n11499), .Y(n17938) );
  OAI22XL U22990 ( .A0(n18541), .A1(n17938), .B0(n18539), .B1(n17901), .Y(
        n17944) );
  XNOR2X1 U22991 ( .A(n18118), .B(n3190), .Y(n17907) );
  OAI22XL U22992 ( .A0(n18107), .A1(n17943), .B0(n18235), .B1(n17907), .Y(
        n17949) );
  XNOR2X1 U22993 ( .A(n18006), .B(n3021), .Y(n17934) );
  ADDFHX1 U22994 ( .A(n17922), .B(n17921), .CI(n17920), .CO(n18369), .S(n17932) );
  ADDFHX1 U22995 ( .A(n17925), .B(n17924), .CI(n17923), .CO(n18352), .S(n17912) );
  ADDFHX1 U22996 ( .A(n17928), .B(n17927), .CI(n17926), .CO(n18367), .S(n18351) );
  CMPR32X1 U22997 ( .A(n17931), .B(n17930), .C(n17929), .CO(n18365), .S(n18350) );
  OAI22X1 U22998 ( .A0(n18226), .A1(n17963), .B0(n17934), .B1(n18223), .Y(
        n17966) );
  XNOR2X1 U22999 ( .A(n18468), .B(M3_mult_x_15_b_1_), .Y(n17968) );
  XNOR2X1 U23000 ( .A(n18503), .B(n3197), .Y(n17967) );
  OAI22XL U23001 ( .A0(n18541), .A1(n17970), .B0(n18539), .B1(n17938), .Y(
        n17976) );
  OAI22X1 U23002 ( .A0(n18239), .A1(n17992), .B0(n18238), .B1(n17941), .Y(
        n17981) );
  XNOR2X1 U23003 ( .A(n18500), .B(n2974), .Y(n17974) );
  OAI22X1 U23004 ( .A0(n18083), .A1(n17974), .B0(n18429), .B1(n17942), .Y(
        n17980) );
  OAI22XL U23005 ( .A0(n18107), .A1(n17975), .B0(n18235), .B1(n17943), .Y(
        n17979) );
  XNOR2X1 U23006 ( .A(n18503), .B(n3049), .Y(n17999) );
  XNOR2X1 U23007 ( .A(n18453), .B(M3_mult_x_15_b_2_), .Y(n17995) );
  OAI22XL U23008 ( .A0(n18541), .A1(n17995), .B0(n18539), .B1(n17970), .Y(
        n18002) );
  XNOR2X1 U23009 ( .A(n3206), .B(n12561), .Y(n18001) );
  OAI22XL U23010 ( .A0(n18242), .A1(n18001), .B0(n18168), .B1(n17973), .Y(
        n18019) );
  XNOR2XL U23011 ( .A(n18500), .B(n11499), .Y(n18000) );
  NOR2BX1 U23012 ( .AN(n2978), .B(n3195), .Y(n18025) );
  XNOR2XL U23013 ( .A(n18006), .B(M3_mult_x_15_b_13_), .Y(n18007) );
  OAI22X1 U23014 ( .A0(n18226), .A1(n18007), .B0(n17994), .B1(n18223), .Y(
        n18024) );
  XNOR2X1 U23015 ( .A(n18500), .B(M3_mult_x_15_b_3_), .Y(n18043) );
  OAI22X1 U23016 ( .A0(n18083), .A1(n18043), .B0(n18429), .B1(n18000), .Y(
        n18030) );
  XNOR2XL U23017 ( .A(n3206), .B(M3_mult_x_15_b_11_), .Y(n18027) );
  OAI22XL U23018 ( .A0(n18242), .A1(n18027), .B0(n18168), .B1(n18001), .Y(
        n18029) );
  ADDFHX1 U23019 ( .A(n18004), .B(n18003), .CI(n18002), .CO(n17996), .S(n18039) );
  OAI22XL U23020 ( .A0(n18239), .A1(n18028), .B0(n18238), .B1(n18005), .Y(
        n18046) );
  XNOR2X1 U23021 ( .A(n18118), .B(n3197), .Y(n18041) );
  XNOR2X1 U23022 ( .A(n18006), .B(n12561), .Y(n18049) );
  OAI22XL U23023 ( .A0(n18177), .A1(n18049), .B0(n18007), .B1(n18223), .Y(
        n18048) );
  OAI22XL U23024 ( .A0(n18541), .A1(n3210), .B0(n5893), .B1(n18008), .Y(n18047) );
  ADDFHX1 U23025 ( .A(n18025), .B(n18024), .CI(n18023), .CO(n18020), .S(n18059) );
  XNOR2XL U23026 ( .A(n3206), .B(M4_mult_x_15_n1680), .Y(n18052) );
  XNOR2X1 U23027 ( .A(n18150), .B(n5430), .Y(n18053) );
  OAI22XL U23028 ( .A0(n18239), .A1(n18053), .B0(n18238), .B1(n18028), .Y(
        n18063) );
  NOR2XL U23029 ( .A(n18314), .B(n18313), .Y(n18035) );
  INVXL U23030 ( .A(n18035), .Y(n18036) );
  NAND2XL U23031 ( .A(n18318), .B(n18036), .Y(n18037) );
  NOR2X1 U23032 ( .A(n18328), .B(n18037), .Y(n18331) );
  XNOR2X1 U23033 ( .A(n18118), .B(n3049), .Y(n18051) );
  OAI22XL U23034 ( .A0(n18107), .A1(n18051), .B0(n18235), .B1(n18041), .Y(
        n18062) );
  OAI22XL U23035 ( .A0(n18083), .A1(n18050), .B0(n18429), .B1(n18043), .Y(
        n18060) );
  CMPR32X1 U23036 ( .A(n18046), .B(n18045), .C(n18044), .CO(n18038), .S(n18073) );
  ADDHXL U23037 ( .A(n18048), .B(n18047), .CO(n18044), .S(n18080) );
  XNOR2X1 U23038 ( .A(n18006), .B(n3190), .Y(n18067) );
  XNOR2X1 U23039 ( .A(n18118), .B(n2974), .Y(n18081) );
  OAI22XL U23040 ( .A0(n18107), .A1(n18081), .B0(n18235), .B1(n18051), .Y(
        n18091) );
  XNOR2XL U23041 ( .A(n3206), .B(M3_mult_x_15_b_9_), .Y(n18084) );
  OAI22X1 U23042 ( .A0(n18242), .A1(n18084), .B0(n18168), .B1(n18052), .Y(
        n18090) );
  XNOR2X1 U23043 ( .A(n18150), .B(n3197), .Y(n18085) );
  OAI22XL U23044 ( .A0(n18239), .A1(n18085), .B0(n18238), .B1(n18053), .Y(
        n18089) );
  ADDFHX1 U23045 ( .A(n18059), .B(n18058), .CI(n18057), .CO(n18054), .S(n18077) );
  OAI22XL U23046 ( .A0(n18111), .A1(n18086), .B0(n18504), .B1(n18066), .Y(
        n18276) );
  NAND2BX1 U23047 ( .AN(n2978), .B(n18500), .Y(n18068) );
  ADDFHX1 U23048 ( .A(n18071), .B(n18069), .CI(n18070), .CO(n18079), .S(n18274) );
  CMPR32X1 U23049 ( .A(n4734), .B(n18079), .C(n18078), .CO(n18072), .S(n18273)
         );
  OAI22XL U23050 ( .A0(n18107), .A1(n18234), .B0(n18235), .B1(n18081), .Y(
        n18245) );
  XNOR2XL U23051 ( .A(n18500), .B(n2978), .Y(n18082) );
  XNOR2X1 U23052 ( .A(n3206), .B(n5430), .Y(n18240) );
  OAI22XL U23053 ( .A0(n18242), .A1(n18240), .B0(n18168), .B1(n18084), .Y(
        n18243) );
  XNOR2X1 U23054 ( .A(n18150), .B(n3049), .Y(n18237) );
  OAI22XL U23055 ( .A0(n18239), .A1(n18237), .B0(n18238), .B1(n18085), .Y(
        n18219) );
  NOR2XL U23056 ( .A(n18300), .B(n18299), .Y(n18095) );
  NOR2XL U23057 ( .A(n18305), .B(n18095), .Y(n18102) );
  NAND2XL U23058 ( .A(n18102), .B(n4620), .Y(n18312) );
  XNOR2X1 U23059 ( .A(n18118), .B(M3_mult_x_15_b_2_), .Y(n18113) );
  OAI22XL U23060 ( .A0(n18107), .A1(n18113), .B0(n18235), .B1(n18236), .Y(
        n18230) );
  XNOR2XL U23061 ( .A(n18503), .B(n2978), .Y(n18103) );
  XNOR2X1 U23062 ( .A(n3206), .B(n2974), .Y(n18117) );
  XNOR2X1 U23063 ( .A(n3206), .B(n3049), .Y(n18108) );
  OAI22XL U23064 ( .A0(n18242), .A1(n18117), .B0(n18168), .B1(n18108), .Y(
        n18123) );
  XNOR2X1 U23065 ( .A(n18150), .B(M3_mult_x_15_b_3_), .Y(n18120) );
  XNOR2X1 U23066 ( .A(n18006), .B(n3049), .Y(n18129) );
  XNOR2X1 U23067 ( .A(n18006), .B(n3197), .Y(n18112) );
  OAI22XL U23068 ( .A0(n18177), .A1(n18129), .B0(n18112), .B1(n18223), .Y(
        n18128) );
  OAI22XL U23069 ( .A0(n18107), .A1(n18106), .B0(n17902), .B1(n18105), .Y(
        n18127) );
  NAND2BX1 U23070 ( .AN(n2978), .B(n18503), .Y(n18109) );
  NOR2BX1 U23071 ( .AN(n2978), .B(n18504), .Y(n18116) );
  OAI22XL U23072 ( .A0(n18242), .A1(n18138), .B0(n18168), .B1(n18117), .Y(
        n18133) );
  XNOR2XL U23073 ( .A(n18118), .B(n2978), .Y(n18119) );
  XNOR2X1 U23074 ( .A(n18150), .B(n12271), .Y(n18130) );
  CMPR32X1 U23075 ( .A(n18123), .B(n18122), .C(n18121), .CO(n18259), .S(n18124) );
  ADDHXL U23076 ( .A(n18128), .B(n18127), .CO(n18121), .S(n18137) );
  NOR2BX1 U23077 ( .AN(n2978), .B(n18235), .Y(n18145) );
  XNOR2X1 U23078 ( .A(n18006), .B(n2974), .Y(n18139) );
  XNOR2X1 U23079 ( .A(n18150), .B(M3_mult_x_15_b_1_), .Y(n18151) );
  OAI22XL U23080 ( .A0(n18239), .A1(n18151), .B0(n18238), .B1(n18130), .Y(
        n18143) );
  CMPR32X1 U23081 ( .A(n18133), .B(n18132), .C(n18131), .CO(n18125), .S(n18135) );
  NOR2XL U23082 ( .A(n18209), .B(n18208), .Y(n18134) );
  ADDFHX1 U23083 ( .A(n18137), .B(n18136), .CI(n18135), .CO(n18208), .S(n18201) );
  OAI22XL U23084 ( .A0(n18177), .A1(n18175), .B0(n18139), .B1(n18223), .Y(
        n18154) );
  NAND2BX1 U23085 ( .AN(n2978), .B(n18150), .Y(n18140) );
  OAI22XL U23086 ( .A0(n18239), .A1(n18152), .B0(n18238), .B1(n18151), .Y(
        n18188) );
  ADDHXL U23087 ( .A(n18154), .B(n18153), .CO(n18147), .S(n18187) );
  OR2X2 U23088 ( .A(n18199), .B(n18198), .Y(n18155) );
  NAND2XL U23089 ( .A(n18204), .B(n18155), .Y(n18207) );
  XNOR2X1 U23090 ( .A(n18006), .B(n12271), .Y(n18165) );
  INVXL U23091 ( .A(n18161), .Y(n18164) );
  INVXL U23092 ( .A(n18157), .Y(n18158) );
  NAND2XL U23093 ( .A(n18159), .B(n18158), .Y(n18163) );
  NAND2XL U23094 ( .A(n18161), .B(n18160), .Y(n18162) );
  OAI21XL U23095 ( .A0(n18164), .A1(n18163), .B0(n18162), .Y(n18174) );
  NAND2BX1 U23096 ( .AN(n2978), .B(n3206), .Y(n18167) );
  NOR2XL U23097 ( .A(n18183), .B(n18182), .Y(n18185) );
  NAND2XL U23098 ( .A(n18183), .B(n18182), .Y(n18184) );
  OAI21XL U23099 ( .A0(n18186), .A1(n18185), .B0(n18184), .Y(n18197) );
  CMPR32X1 U23100 ( .A(n18189), .B(n18188), .C(n18187), .CO(n18198), .S(n18195) );
  CMPR32X1 U23101 ( .A(n18192), .B(n18191), .C(n18190), .CO(n18194), .S(n18183) );
  AND2X2 U23102 ( .A(n18195), .B(n18194), .Y(n18196) );
  AOI21XL U23103 ( .A0(n18197), .A1(n18193), .B0(n18196), .Y(n18206) );
  AND2X2 U23104 ( .A(n18201), .B(n18200), .Y(n18202) );
  AOI21XL U23105 ( .A0(n18204), .A1(n18203), .B0(n18202), .Y(n18205) );
  OAI21XL U23106 ( .A0(n18207), .A1(n18206), .B0(n18205), .Y(n18215) );
  NAND2XL U23107 ( .A(n18209), .B(n18208), .Y(n18213) );
  NAND2XL U23108 ( .A(n18211), .B(n18210), .Y(n18212) );
  AOI21XL U23109 ( .A0(n18216), .A1(n18215), .B0(n18214), .Y(n18270) );
  CMPR32X1 U23110 ( .A(n18219), .B(n18218), .C(n18217), .CO(n18281), .S(n18288) );
  OAI22X1 U23111 ( .A0(n18226), .A1(n18225), .B0(n18224), .B1(n18223), .Y(
        n18232) );
  ADDFHX1 U23112 ( .A(n18230), .B(n18229), .CI(n18228), .CO(n18252), .S(n18260) );
  OAI22XL U23113 ( .A0(n18242), .A1(n18241), .B0(n18168), .B1(n18240), .Y(
        n18246) );
  CMPR32X1 U23114 ( .A(n18245), .B(n18244), .C(n18243), .CO(n18282), .S(n18277) );
  CMPR32X1 U23115 ( .A(n18248), .B(n18247), .C(n18246), .CO(n18278), .S(n18257) );
  ADDFHX1 U23116 ( .A(n18257), .B(n18256), .CI(n18255), .CO(n18264), .S(n18263) );
  OR2X2 U23117 ( .A(n18263), .B(n18262), .Y(n18261) );
  AND2X2 U23118 ( .A(n18263), .B(n18262), .Y(n18266) );
  OAI21XL U23119 ( .A0(n18270), .A1(n18269), .B0(n18268), .Y(n18298) );
  NOR2XL U23120 ( .A(n18291), .B(n18290), .Y(n18289) );
  NOR2XL U23121 ( .A(n18295), .B(n18289), .Y(n18297) );
  NAND2XL U23122 ( .A(n18291), .B(n18290), .Y(n18294) );
  AND2X2 U23123 ( .A(n18307), .B(n18306), .Y(n18308) );
  AOI21X1 U23124 ( .A0(n18309), .A1(n4620), .B0(n18308), .Y(n18310) );
  OAI21X1 U23125 ( .A0(n18312), .A1(n18311), .B0(n18310), .Y(n18330) );
  CMPR32X1 U23126 ( .A(n18346), .B(n18345), .C(n18344), .CO(n18341), .S(n18376) );
  ADDFHX4 U23127 ( .A(n18355), .B(n18354), .CI(n18353), .CO(n18333), .S(n18356) );
  ADDFHX1 U23128 ( .A(n18370), .B(n18369), .CI(n18368), .CO(n18380), .S(n18385) );
  OAI21XL U23129 ( .A0(n18881), .A1(n18875), .B0(n18882), .Y(n18418) );
  AOI21X1 U23130 ( .A0(n18867), .A1(n18419), .B0(n18418), .Y(n18420) );
  XNOR2X1 U23131 ( .A(M4_a_17_), .B(n3196), .Y(n18432) );
  XNOR2X1 U23132 ( .A(n18604), .B(n3048), .Y(n18425) );
  OAI22XL U23133 ( .A0(n18624), .A1(n18432), .B0(n18625), .B1(n18425), .Y(
        n18437) );
  XNOR2X1 U23134 ( .A(n18453), .B(n3202), .Y(n18433) );
  XNOR2XL U23135 ( .A(n18468), .B(M3_mult_x_15_b_21_), .Y(n18424) );
  OAI22XL U23136 ( .A0(n18522), .A1(n18434), .B0(n3195), .B1(n18424), .Y(
        n18440) );
  XNOR2X1 U23137 ( .A(n25883), .B(n18611), .Y(n18431) );
  XNOR2X1 U23138 ( .A(n25883), .B(n3198), .Y(n18426) );
  OAI22XL U23139 ( .A0(n18659), .A1(n18431), .B0(n17832), .B1(n18426), .Y(
        n18439) );
  XNOR2X1 U23140 ( .A(n18638), .B(n3021), .Y(n18430) );
  XNOR2X1 U23141 ( .A(n18638), .B(n3201), .Y(n18423) );
  OAI22XL U23142 ( .A0(n18652), .A1(n18430), .B0(n18653), .B1(n18423), .Y(
        n18438) );
  XNOR2X1 U23143 ( .A(n18638), .B(n3196), .Y(n18451) );
  OAI22XL U23144 ( .A0(n18652), .A1(n18423), .B0(n18653), .B1(n18451), .Y(
        n18450) );
  XNOR2X1 U23145 ( .A(n18468), .B(n3202), .Y(n18452) );
  OAI22XL U23146 ( .A0(n18522), .A1(n18424), .B0(n3195), .B1(n18452), .Y(
        n18449) );
  OAI22XL U23147 ( .A0(n18624), .A1(n18425), .B0(n18625), .B1(n18444), .Y(
        n18448) );
  XNOR2X1 U23148 ( .A(n25883), .B(n3021), .Y(n18445) );
  OAI22XL U23149 ( .A0(n18666), .A1(n18426), .B0(n17832), .B1(n18445), .Y(
        n18443) );
  OAI22XL U23150 ( .A0(n18721), .A1(n12561), .B0(n17512), .B1(
        M3_mult_x_15_b_13_), .Y(n18427) );
  OAI22XL U23151 ( .A0(n18541), .A1(n18453), .B0(n18539), .B1(n3210), .Y(
        n18446) );
  OAI22X1 U23152 ( .A0(n18721), .A1(n3190), .B0(n17512), .B1(n12561), .Y(
        n18497) );
  OAI22XL U23153 ( .A0(n18083), .A1(n18500), .B0(n18429), .B1(n18428), .Y(
        n18496) );
  OAI22XL U23154 ( .A0(n18652), .A1(n18544), .B0(n18653), .B1(n18430), .Y(
        n18507) );
  XNOR2XL U23155 ( .A(n25883), .B(M3_mult_x_15_b_13_), .Y(n18542) );
  OAI22XL U23156 ( .A0(n18624), .A1(n18499), .B0(n18625), .B1(n18432), .Y(
        n18505) );
  XNOR2XL U23157 ( .A(n18453), .B(M3_mult_x_15_b_21_), .Y(n18538) );
  OAI22XL U23158 ( .A0(n18721), .A1(M4_mult_x_15_n1680), .B0(n17512), .B1(
        n3190), .Y(n18523) );
  CMPR32X1 U23159 ( .A(n18437), .B(n18436), .C(n18435), .CO(n18492), .S(n18509) );
  CMPR32X1 U23160 ( .A(n18440), .B(n18439), .C(n18438), .CO(n18491), .S(n18508) );
  XNOR2X1 U23161 ( .A(M4_a_17_), .B(M3_mult_x_15_b_21_), .Y(n18462) );
  OAI22XL U23162 ( .A0(n18624), .A1(n18444), .B0(n18625), .B1(n18462), .Y(
        n18465) );
  XNOR2X1 U23163 ( .A(n25883), .B(n3201), .Y(n18460) );
  OAI22XL U23164 ( .A0(n18666), .A1(n18445), .B0(n17832), .B1(n18460), .Y(
        n18464) );
  OAI22XL U23165 ( .A0(n18721), .A1(n18611), .B0(n17512), .B1(n3198), .Y(
        n18466) );
  CMPR32X1 U23166 ( .A(n18450), .B(n18449), .C(n18448), .CO(n18455), .S(n18490) );
  OAI22XL U23167 ( .A0(n18652), .A1(n18451), .B0(n18653), .B1(n18461), .Y(
        n18471) );
  XNOR2X1 U23168 ( .A(n25883), .B(n3196), .Y(n18482) );
  OAI22XL U23169 ( .A0(n18666), .A1(n18460), .B0(n17832), .B1(n18482), .Y(
        n18480) );
  XNOR2X1 U23170 ( .A(n18604), .B(n3202), .Y(n18484) );
  CMPR32X1 U23171 ( .A(n18465), .B(n18464), .C(n18463), .CO(n18488), .S(n18458) );
  CMPR32X1 U23172 ( .A(n12561), .B(n12518), .C(n18466), .CO(n18477), .S(n18463) );
  NOR2X1 U23173 ( .A(n18686), .B(n18685), .Y(n18941) );
  XNOR2XL U23174 ( .A(n18638), .B(M3_mult_x_15_b_21_), .Y(n18608) );
  OAI22XL U23175 ( .A0(n18652), .A1(n18481), .B0(n18653), .B1(n18608), .Y(
        n18607) );
  XNOR2X1 U23176 ( .A(n25883), .B(n3048), .Y(n18609) );
  OAI22XL U23177 ( .A0(n18721), .A1(n3021), .B0(n17512), .B1(n3201), .Y(n18610) );
  CMPR32X1 U23178 ( .A(n18489), .B(n18488), .C(n18487), .CO(n18597), .S(n18472) );
  CMPR32X1 U23179 ( .A(n18492), .B(n18491), .C(n18490), .CO(n18516), .S(n18574) );
  OAI22XL U23180 ( .A0(n18083), .A1(n18502), .B0(n18501), .B1(n18500), .Y(
        n18536) );
  OAI2BB1XL U23181 ( .A0N(n18504), .A1N(n18111), .B0(n18503), .Y(n18535) );
  CMPR32X1 U23182 ( .A(n18513), .B(n18512), .C(n18511), .CO(n18515), .S(n18572) );
  OAI22XL U23183 ( .A0(n18522), .A1(n18521), .B0(n3195), .B1(n18520), .Y(
        n18553) );
  CMPR32X1 U23184 ( .A(n18537), .B(n18536), .C(n18535), .CO(n18530), .S(n18558) );
  OAI22XL U23185 ( .A0(n18541), .A1(n18540), .B0(n18539), .B1(n18538), .Y(
        n18548) );
  CMPR32X1 U23186 ( .A(n18556), .B(n18555), .C(n18554), .CO(n18587), .S(n18589) );
  CMPR32X1 U23187 ( .A(n18562), .B(n18561), .C(n18560), .CO(n18596), .S(n18585) );
  NOR2X1 U23188 ( .A(n18681), .B(n18680), .Y(n18578) );
  INVX1 U23189 ( .A(n18578), .Y(n18855) );
  NOR2X2 U23190 ( .A(n18692), .B(n18926), .Y(n18694) );
  ADDFHX1 U23191 ( .A(n18584), .B(n18583), .CI(n18582), .CO(n18593), .S(n18588) );
  NOR2X1 U23192 ( .A(n18861), .B(n18857), .Y(n18846) );
  OAI22XL U23193 ( .A0(n18721), .A1(n3201), .B0(n17512), .B1(n3196), .Y(n18622) );
  OAI22XL U23194 ( .A0(n18652), .A1(n18608), .B0(n18653), .B1(n18623), .Y(
        n18620) );
  CMPR32X1 U23195 ( .A(n18611), .B(n3198), .C(n18610), .CO(n18618), .S(n18601)
         );
  CMPR32X1 U23196 ( .A(n18614), .B(n18613), .C(n18612), .CO(n18615), .S(n18598) );
  CMPR32X1 U23197 ( .A(n18617), .B(n18616), .C(n18615), .CO(n18698), .S(n18695) );
  CMPR32X1 U23198 ( .A(n18620), .B(n18619), .C(n18618), .CO(n18631), .S(n18626) );
  OAI22XL U23199 ( .A0(n18721), .A1(n3196), .B0(n17512), .B1(n3048), .Y(n18636) );
  CMPR32X1 U23200 ( .A(n3043), .B(n18622), .C(n18621), .CO(n18641), .S(n18628)
         );
  OAI2BB1XL U23201 ( .A0N(n18625), .A1N(n18624), .B0(M4_a_17_), .Y(n18632) );
  CMPR32X1 U23202 ( .A(n18634), .B(n18633), .C(n18632), .CO(n18645), .S(n18640) );
  CMPR32X1 U23203 ( .A(n3021), .B(n3201), .C(n18636), .CO(n18649), .S(n18642)
         );
  CMPR32X1 U23204 ( .A(n18645), .B(n18644), .C(n18643), .CO(n18705), .S(n18699) );
  CMPR32X1 U23205 ( .A(n18650), .B(n18649), .C(n18648), .CO(n18655), .S(n18644) );
  CMPR32X1 U23206 ( .A(n18656), .B(n18655), .C(n18654), .CO(n18707), .S(n18704) );
  CMPR32X1 U23207 ( .A(n3196), .B(n3048), .C(n18657), .CO(n18665), .S(n18660)
         );
  CMPR32X1 U23208 ( .A(n18662), .B(n18661), .C(n18660), .CO(n18663), .S(n18654) );
  CMPR32X1 U23209 ( .A(n18665), .B(n18664), .C(n18663), .CO(n18711), .S(n18706) );
  CMPR32X1 U23210 ( .A(n5960), .B(n18668), .C(n18667), .CO(n18669), .S(n18664)
         );
  CMPR32X1 U23211 ( .A(n18671), .B(n18670), .C(n18669), .CO(n18713), .S(n18710) );
  CMPR32X1 U23212 ( .A(n18673), .B(M3_mult_x_15_b_21_), .C(n18672), .CO(n18720), .S(n18670) );
  OR2X2 U23213 ( .A(n18713), .B(n18712), .Y(n18997) );
  NAND2X1 U23214 ( .A(n18679), .B(n18678), .Y(n18848) );
  NAND2XL U23215 ( .A(n18681), .B(n18680), .Y(n18854) );
  INVXL U23216 ( .A(n18854), .Y(n18682) );
  NAND2XL U23217 ( .A(n18684), .B(n18683), .Y(n18931) );
  INVXL U23218 ( .A(n18931), .Y(n18934) );
  NAND2XL U23219 ( .A(n18688), .B(n18687), .Y(n18952) );
  OAI21XL U23220 ( .A0(n18951), .A1(n18945), .B0(n18952), .Y(n18689) );
  AOI21XL U23221 ( .A0(n18961), .A1(n18966), .B0(n18701), .Y(n18702) );
  OAI21XL U23222 ( .A0(n18988), .A1(n19003), .B0(n18989), .Y(n18708) );
  CMPR32X1 U23223 ( .A(n5957), .B(n4227), .C(n18720), .CO(n18724), .S(n18712)
         );
  INVXL U23224 ( .A(n18727), .Y(n18730) );
  INVXL U23225 ( .A(n18728), .Y(n18729) );
  AOI21XL U23226 ( .A0(n18792), .A1(n18730), .B0(n18729), .Y(n18735) );
  INVXL U23227 ( .A(n18731), .Y(n18733) );
  NAND2XL U23228 ( .A(n18733), .B(n18732), .Y(n18734) );
  OAI21XL U23229 ( .A0(n26304), .A1(n17167), .B0(n18736), .Y(n18738) );
  OAI21XL U23230 ( .A0(n26285), .A1(n17167), .B0(n18739), .Y(n18740) );
  OAI21XL U23231 ( .A0(n26284), .A1(n15940), .B0(n18741), .Y(n18743) );
  AND2X2 U23232 ( .A(n3111), .B(data[88]), .Y(n18742) );
  NOR2X1 U23233 ( .A(n18743), .B(n18742), .Y(n19027) );
  OAI21XL U23234 ( .A0(n26298), .A1(n17167), .B0(n18747), .Y(n18749) );
  OAI21XL U23235 ( .A0(n26044), .A1(n15940), .B0(n18753), .Y(n18755) );
  CMPR32X1 U23236 ( .A(n18770), .B(n18769), .C(n18768), .CO(n18765), .S(n25124) );
  CMPR32X1 U23237 ( .A(n18773), .B(n18772), .C(n18771), .CO(n18784), .S(n20795) );
  CMPR32X1 U23238 ( .A(n18776), .B(n18775), .C(n18774), .CO(n18771), .S(n24348) );
  CMPR32X1 U23239 ( .A(n18779), .B(n18778), .C(n18777), .CO(n18774), .S(n20787) );
  CMPR22X1 U23240 ( .A(n19026), .B(n18780), .CO(n18777), .S(n20786) );
  CMPR32X1 U23241 ( .A(n18783), .B(n18782), .C(n18781), .CO(n18768), .S(n24110) );
  CMPR32X1 U23242 ( .A(n18786), .B(n18785), .C(n18784), .CO(n18781), .S(n24275) );
  NAND4BXL U23243 ( .AN(n25124), .B(n18789), .C(n18788), .D(n18787), .Y(n18790) );
  NOR3X1 U23244 ( .A(n20649), .B(n25129), .C(n18790), .Y(n18968) );
  INVXL U23245 ( .A(n18968), .Y(n18829) );
  INVXL U23246 ( .A(n18832), .Y(n18793) );
  OAI21XL U23247 ( .A0(n18817), .A1(n18818), .B0(n18820), .Y(n18796) );
  OAI21XL U23248 ( .A0(n18797), .A1(M4_U3_U1_enc_tree_2__4__16_), .B0(n18796), 
        .Y(n18802) );
  OAI21X1 U23249 ( .A0(n18833), .A1(n18832), .B0(n18831), .Y(n18838) );
  XNOR2X2 U23250 ( .A(n18838), .B(n18837), .Y(n18973) );
  OAI21XL U23251 ( .A0(n18973), .A1(n18844), .B0(n24250), .Y(n18845) );
  INVXL U23252 ( .A(n18846), .Y(n18933) );
  OAI21X2 U23253 ( .A0(n19014), .A1(n18933), .B0(n18938), .Y(n18850) );
  NAND2XL U23254 ( .A(n18846), .B(n18847), .Y(n18853) );
  INVXL U23255 ( .A(n18857), .Y(n18859) );
  INVXL U23256 ( .A(n18861), .Y(n18863) );
  INVXL U23257 ( .A(n18865), .Y(n18874) );
  NAND2XL U23258 ( .A(n18895), .B(n18865), .Y(n18869) );
  INVXL U23259 ( .A(n18867), .Y(n18876) );
  NAND2XL U23260 ( .A(n18873), .B(n18875), .Y(n18871) );
  NOR2XL U23261 ( .A(n18874), .B(n18870), .Y(n18878) );
  NAND2XL U23262 ( .A(n18878), .B(n18895), .Y(n18880) );
  OAI21XL U23263 ( .A0(n18876), .A1(n18870), .B0(n18875), .Y(n18877) );
  AOI21XL U23264 ( .A0(n18878), .A1(n18896), .B0(n18877), .Y(n18879) );
  INVXL U23265 ( .A(n18881), .Y(n18883) );
  NAND2XL U23266 ( .A(n18883), .B(n18882), .Y(n18884) );
  XNOR2X2 U23267 ( .A(n18885), .B(n18884), .Y(n23515) );
  NAND2XL U23268 ( .A(n18895), .B(n18900), .Y(n18889) );
  INVXL U23269 ( .A(n18899), .Y(n18887) );
  INVXL U23270 ( .A(n18890), .Y(n18892) );
  NAND2XL U23271 ( .A(n18892), .B(n18891), .Y(n18893) );
  XNOR2X1 U23272 ( .A(n18894), .B(n18893), .Y(n23529) );
  INVXL U23273 ( .A(n18895), .Y(n18898) );
  INVXL U23274 ( .A(n18896), .Y(n18897) );
  OAI21X1 U23275 ( .A0(n18925), .A1(n18898), .B0(n18897), .Y(n18902) );
  INVXL U23276 ( .A(n18903), .Y(n18906) );
  INVXL U23277 ( .A(n18904), .Y(n18905) );
  INVXL U23278 ( .A(n18907), .Y(n18911) );
  NAND2XL U23279 ( .A(n18903), .B(n18911), .Y(n18913) );
  INVXL U23280 ( .A(n18909), .Y(n18910) );
  AOI21XL U23281 ( .A0(n18904), .A1(n18911), .B0(n18910), .Y(n18912) );
  INVXL U23282 ( .A(n18923), .Y(n18917) );
  INVXL U23283 ( .A(n18919), .Y(n18921) );
  INVXL U23284 ( .A(n18926), .Y(n18932) );
  NAND2XL U23285 ( .A(n18846), .B(n18932), .Y(n18930) );
  INVXL U23286 ( .A(n18927), .Y(n18935) );
  NAND2XL U23287 ( .A(n18932), .B(n3000), .Y(n18937) );
  NOR2XL U23288 ( .A(n18933), .B(n18937), .Y(n18944) );
  INVXL U23289 ( .A(n18944), .Y(n18940) );
  OAI21XL U23290 ( .A0(n18938), .A1(n18937), .B0(n18936), .Y(n18948) );
  INVXL U23291 ( .A(n18984), .Y(n19011) );
  NAND2XL U23292 ( .A(n18944), .B(n18947), .Y(n18950) );
  INVXL U23293 ( .A(n18945), .Y(n18946) );
  INVXL U23294 ( .A(n18951), .Y(n18953) );
  INVXL U23295 ( .A(n18960), .Y(n18958) );
  OAI21X1 U23296 ( .A0(n18984), .A1(n18942), .B0(n18956), .Y(n18963) );
  NAND2XL U23297 ( .A(n18960), .B(n18962), .Y(n18965) );
  NOR3X1 U23298 ( .A(n18968), .B(n20649), .C(n18970), .Y(n19023) );
  NAND3X1 U23299 ( .A(n23513), .B(n23529), .C(n18972), .Y(n18977) );
  NAND4BX2 U23300 ( .AN(n18974), .B(n23454), .C(n23460), .D(n23458), .Y(n18976) );
  INVXL U23301 ( .A(n18979), .Y(n18983) );
  NAND2XL U23302 ( .A(n18999), .B(n19004), .Y(n18987) );
  OAI21XL U23303 ( .A0(n18984), .A1(n18983), .B0(n18982), .Y(n19000) );
  AOI21XL U23304 ( .A0(n19000), .A1(n19004), .B0(n18985), .Y(n18986) );
  OAI21X1 U23305 ( .A0(n19014), .A1(n18987), .B0(n18986), .Y(n18991) );
  NAND2XL U23306 ( .A(n19007), .B(n18992), .Y(n18995) );
  AOI21XL U23307 ( .A0(n19011), .A1(n18992), .B0(n18993), .Y(n18994) );
  INVXL U23308 ( .A(n19006), .Y(n19010) );
  NAND2XL U23309 ( .A(n19007), .B(n19010), .Y(n19013) );
  NAND2X1 U23310 ( .A(n22482), .B(n22481), .Y(n20653) );
  AOI22XL U23311 ( .A0(n24244), .A1(n25636), .B0(n2983), .B1(temp2[18]), .Y(
        n19046) );
  NAND2XL U23312 ( .A(n24236), .B(n25638), .Y(n19045) );
  NOR2XL U23313 ( .A(n5033), .B(n19050), .Y(n19049) );
  AOI22XL U23314 ( .A0(n24210), .A1(n25636), .B0(n2984), .B1(temp2[14]), .Y(
        n19052) );
  NAND2XL U23315 ( .A(n24199), .B(n25638), .Y(n19051) );
  INVXL U23316 ( .A(n19053), .Y(n19055) );
  NAND2XL U23317 ( .A(n19055), .B(n19054), .Y(n19056) );
  XOR2X1 U23318 ( .A(n19056), .B(n20947), .Y(n20950) );
  XNOR2X1 U23319 ( .A(n23738), .B(n19057), .Y(n19075) );
  XNOR2X1 U23320 ( .A(n5100), .B(n19058), .Y(n19079) );
  INVXL U23321 ( .A(n19059), .Y(n19061) );
  NAND2XL U23322 ( .A(n19061), .B(n19060), .Y(n19062) );
  AOI22XL U23323 ( .A0(n23949), .A1(n19083), .B0(n23947), .B1(n20962), .Y(
        n19068) );
  NAND2XL U23324 ( .A(n5100), .B(n19076), .Y(n19078) );
  AOI22XL U23325 ( .A0(n23949), .A1(n23725), .B0(n23947), .B1(n19083), .Y(
        n19084) );
  NAND2XL U23326 ( .A(n3141), .B(n19090), .Y(n19094) );
  NOR2XL U23327 ( .A(n19094), .B(n19096), .Y(n19091) );
  INVXL U23328 ( .A(n19094), .Y(n19095) );
  NAND2XL U23329 ( .A(n23744), .B(n19095), .Y(n19097) );
  XOR2X1 U23330 ( .A(n19096), .B(n19097), .Y(n23435) );
  AOI22X1 U23331 ( .A0(n3081), .A1(n23650), .B0(n23435), .B1(n4267), .Y(n24177) );
  INVXL U23332 ( .A(n24177), .Y(n20268) );
  INVXL U23333 ( .A(n19100), .Y(n19101) );
  NAND2X1 U23334 ( .A(n3132), .B(n19101), .Y(n19102) );
  INVXL U23335 ( .A(n19322), .Y(n19107) );
  NAND2X1 U23336 ( .A(n19107), .B(n19278), .Y(n24300) );
  AOI22XL U23337 ( .A0(n3027), .A1(w2[35]), .B0(n19161), .B1(w1[67]), .Y(
        n19108) );
  OAI21XL U23338 ( .A0(n19237), .A1(n25953), .B0(n19108), .Y(n19563) );
  AOI22XL U23339 ( .A0(n19346), .A1(y11[3]), .B0(n19161), .B1(temp2[3]), .Y(
        n19109) );
  OAI21XL U23340 ( .A0(n19237), .A1(n26567), .B0(n19109), .Y(n19562) );
  NOR2XL U23341 ( .A(n19736), .B(n19562), .Y(n19122) );
  AOI22XL U23342 ( .A0(n3027), .A1(w2[34]), .B0(n19161), .B1(w1[66]), .Y(
        n19110) );
  OAI21XL U23343 ( .A0(n19237), .A1(n25954), .B0(n19110), .Y(n19561) );
  AOI22XL U23344 ( .A0(n3027), .A1(y11[2]), .B0(n19161), .B1(temp2[2]), .Y(
        n19111) );
  OAI21XL U23345 ( .A0(n3063), .A1(n26568), .B0(n19111), .Y(n19560) );
  NOR2XL U23346 ( .A(n19720), .B(n19560), .Y(n19112) );
  NOR2XL U23347 ( .A(n19122), .B(n19112), .Y(n19125) );
  AOI22XL U23348 ( .A0(n19349), .A1(w2[33]), .B0(n3026), .B1(w1[65]), .Y(
        n19113) );
  OAI21XL U23349 ( .A0(n19237), .A1(n25955), .B0(n19113), .Y(n19557) );
  AOI22XL U23350 ( .A0(n3027), .A1(y11[1]), .B0(n19161), .B1(temp2[1]), .Y(
        n19114) );
  OAI21XL U23351 ( .A0(n19237), .A1(n26569), .B0(n19114), .Y(n19556) );
  NOR2XL U23352 ( .A(n19598), .B(n19556), .Y(n19119) );
  AOI22XL U23353 ( .A0(n19349), .A1(w2[32]), .B0(n3062), .B1(w1[64]), .Y(
        n19115) );
  OAI21XL U23354 ( .A0(n19237), .A1(n25956), .B0(n19115), .Y(n19555) );
  AOI22XL U23355 ( .A0(n19346), .A1(y11[0]), .B0(n19161), .B1(temp2[0]), .Y(
        n19116) );
  OAI21XL U23356 ( .A0(n3063), .A1(n26570), .B0(n19116), .Y(n19554) );
  NAND2XL U23357 ( .A(n19598), .B(n19556), .Y(n19117) );
  NAND2XL U23358 ( .A(n19720), .B(n19560), .Y(n19121) );
  NAND2XL U23359 ( .A(n19736), .B(n19562), .Y(n19120) );
  OAI21XL U23360 ( .A0(n19122), .A1(n19121), .B0(n19120), .Y(n19123) );
  AOI21XL U23361 ( .A0(n19125), .A1(n19124), .B0(n19123), .Y(n19148) );
  AOI22XL U23362 ( .A0(n3027), .A1(w2[36]), .B0(n19161), .B1(w1[68]), .Y(
        n19126) );
  OAI21XL U23363 ( .A0(n19237), .A1(n25952), .B0(n19126), .Y(n19568) );
  AOI22XL U23364 ( .A0(n19346), .A1(y11[4]), .B0(n19161), .B1(temp2[4]), .Y(
        n19127) );
  OAI21XL U23365 ( .A0(n3063), .A1(n26566), .B0(n19127), .Y(n19567) );
  NOR2XL U23366 ( .A(n19752), .B(n19567), .Y(n19130) );
  AOI22XL U23367 ( .A0(n3027), .A1(w2[37]), .B0(n19161), .B1(w1[69]), .Y(
        n19128) );
  OAI21XL U23368 ( .A0(n19237), .A1(n25951), .B0(n19128), .Y(n19538) );
  AOI22XL U23369 ( .A0(n19346), .A1(y11[5]), .B0(n19161), .B1(temp2[5]), .Y(
        n19129) );
  OAI21XL U23370 ( .A0(n3063), .A1(n26565), .B0(n19129), .Y(n19537) );
  NOR2XL U23371 ( .A(n19130), .B(n19139), .Y(n19136) );
  AOI22XL U23372 ( .A0(n19349), .A1(w2[38]), .B0(n19161), .B1(w1[70]), .Y(
        n19131) );
  OAI21XL U23373 ( .A0(n19237), .A1(n25950), .B0(n19131), .Y(n19485) );
  AOI22XL U23374 ( .A0(n19346), .A1(y11[6]), .B0(n19161), .B1(temp2[6]), .Y(
        n19132) );
  OAI21XL U23375 ( .A0(n3063), .A1(n26564), .B0(n19132), .Y(n19484) );
  NOR2XL U23376 ( .A(n19508), .B(n19484), .Y(n19135) );
  AOI22XL U23377 ( .A0(n3027), .A1(w2[39]), .B0(n19161), .B1(w1[71]), .Y(
        n19133) );
  OAI21XL U23378 ( .A0(n19237), .A1(n25892), .B0(n19133), .Y(n19487) );
  AOI22XL U23379 ( .A0(n19346), .A1(y11[7]), .B0(n19161), .B1(temp2[7]), .Y(
        n19134) );
  OAI21XL U23380 ( .A0(n3063), .A1(n26563), .B0(n19134), .Y(n19486) );
  NOR2X1 U23381 ( .A(n19135), .B(n19142), .Y(n19145) );
  NAND2XL U23382 ( .A(n19136), .B(n19145), .Y(n19147) );
  NAND2XL U23383 ( .A(n19752), .B(n19567), .Y(n19138) );
  NAND2XL U23384 ( .A(n19551), .B(n19537), .Y(n19137) );
  OAI21XL U23385 ( .A0(n19139), .A1(n19138), .B0(n19137), .Y(n19144) );
  NAND2XL U23386 ( .A(n19508), .B(n19484), .Y(n19141) );
  NAND2XL U23387 ( .A(n19532), .B(n19486), .Y(n19140) );
  OAI21XL U23388 ( .A0(n19142), .A1(n19141), .B0(n19140), .Y(n19143) );
  AOI22XL U23389 ( .A0(n3027), .A1(w2[40]), .B0(n19161), .B1(w1[72]), .Y(
        n19149) );
  OAI21XL U23390 ( .A0(n19237), .A1(n25949), .B0(n19149), .Y(n19384) );
  AOI22XL U23391 ( .A0(n19346), .A1(y11[8]), .B0(n19161), .B1(temp2[8]), .Y(
        n19150) );
  OAI21XL U23392 ( .A0(n3063), .A1(n26562), .B0(n19150), .Y(n19383) );
  NOR2XL U23393 ( .A(n19455), .B(n19383), .Y(n19153) );
  AOI22XL U23394 ( .A0(n3027), .A1(w2[41]), .B0(n19161), .B1(w1[73]), .Y(
        n19151) );
  OAI21XL U23395 ( .A0(n19237), .A1(n25891), .B0(n19151), .Y(n19386) );
  AOI22XL U23396 ( .A0(n19346), .A1(y11[9]), .B0(n19161), .B1(temp2[9]), .Y(
        n19152) );
  OAI21XL U23397 ( .A0(n19237), .A1(n26561), .B0(n19152), .Y(n19385) );
  NOR2XL U23398 ( .A(n19153), .B(n19175), .Y(n19159) );
  AOI22XL U23399 ( .A0(n3027), .A1(w2[43]), .B0(n19161), .B1(w1[75]), .Y(
        n19154) );
  OAI21XL U23400 ( .A0(n19237), .A1(n25947), .B0(n19154), .Y(n19393) );
  AOI22XL U23401 ( .A0(n3027), .A1(y11[11]), .B0(n19161), .B1(temp2[11]), .Y(
        n19155) );
  OAI21XL U23402 ( .A0(n3063), .A1(n26559), .B0(n19155), .Y(n19392) );
  AOI22XL U23403 ( .A0(n3027), .A1(w2[42]), .B0(n19161), .B1(w1[74]), .Y(
        n19156) );
  OAI21XL U23404 ( .A0(n19237), .A1(n25948), .B0(n19156), .Y(n19390) );
  AOI22XL U23405 ( .A0(n19346), .A1(y11[10]), .B0(n19161), .B1(temp2[10]), .Y(
        n19157) );
  OAI21XL U23406 ( .A0(n3063), .A1(n26560), .B0(n19157), .Y(n19389) );
  NOR2XL U23407 ( .A(n19787), .B(n19389), .Y(n19158) );
  NAND2XL U23408 ( .A(n19159), .B(n19181), .Y(n19172) );
  AOI22XL U23409 ( .A0(n3027), .A1(w2[44]), .B0(n19161), .B1(w1[76]), .Y(
        n19160) );
  OAI21XL U23410 ( .A0(n19237), .A1(n25946), .B0(n19160), .Y(n19365) );
  AOI22XL U23411 ( .A0(n19346), .A1(y11[12]), .B0(n19161), .B1(temp2[12]), .Y(
        n19162) );
  OAI21XL U23412 ( .A0(n3063), .A1(n26558), .B0(n19162), .Y(n19364) );
  AOI22XL U23413 ( .A0(n19349), .A1(w2[45]), .B0(n19161), .B1(w1[77]), .Y(
        n19163) );
  OAI21XL U23414 ( .A0(n19237), .A1(n25945), .B0(n19163), .Y(n19367) );
  AOI22XL U23415 ( .A0(n3027), .A1(y11[13]), .B0(n19216), .B1(temp2[13]), .Y(
        n19164) );
  OAI21XL U23416 ( .A0(n3063), .A1(n26557), .B0(n19164), .Y(n19366) );
  AOI22XL U23417 ( .A0(n19235), .A1(w2[47]), .B0(n19161), .B1(w1[79]), .Y(
        n19166) );
  OAI21XL U23418 ( .A0(n19237), .A1(n25943), .B0(n19166), .Y(n19374) );
  AOI22XL U23419 ( .A0(n19235), .A1(y11[15]), .B0(n3062), .B1(temp2[15]), .Y(
        n19167) );
  OAI21XL U23420 ( .A0(n3063), .A1(n26555), .B0(n19167), .Y(n19373) );
  AOI22XL U23421 ( .A0(n19235), .A1(w2[46]), .B0(n19161), .B1(w1[78]), .Y(
        n19168) );
  OAI21XL U23422 ( .A0(n3063), .A1(n25944), .B0(n19168), .Y(n19371) );
  AOI22XL U23423 ( .A0(n3027), .A1(y11[14]), .B0(n3026), .B1(temp2[14]), .Y(
        n19169) );
  OAI21XL U23424 ( .A0(n3063), .A1(n26556), .B0(n19169), .Y(n19370) );
  NAND2XL U23425 ( .A(n19479), .B(n19385), .Y(n19173) );
  OAI21XL U23426 ( .A0(n19175), .A1(n19174), .B0(n19173), .Y(n19180) );
  NAND2XL U23427 ( .A(n19787), .B(n19389), .Y(n19177) );
  NAND2XL U23428 ( .A(n19794), .B(n19392), .Y(n19176) );
  OAI21XL U23429 ( .A0(n19178), .A1(n19177), .B0(n19176), .Y(n19179) );
  AOI21XL U23430 ( .A0(n19181), .A1(n19180), .B0(n19179), .Y(n19193) );
  NAND2XL U23431 ( .A(n19802), .B(n19364), .Y(n19183) );
  NAND2XL U23432 ( .A(n19810), .B(n19366), .Y(n19182) );
  OAI21XL U23433 ( .A0(n19184), .A1(n19183), .B0(n19182), .Y(n19189) );
  NAND2XL U23434 ( .A(n19815), .B(n19370), .Y(n19186) );
  NAND2XL U23435 ( .A(n19820), .B(n19373), .Y(n19185) );
  OAI21XL U23436 ( .A0(n19187), .A1(n19186), .B0(n19185), .Y(n19188) );
  AOI21X1 U23437 ( .A0(n19196), .A1(n19195), .B0(n19194), .Y(n19289) );
  AOI22XL U23438 ( .A0(n3027), .A1(w2[48]), .B0(n19161), .B1(w1[80]), .Y(
        n19197) );
  OAI21XL U23439 ( .A0(n19237), .A1(n25942), .B0(n19197), .Y(n19436) );
  AOI22XL U23440 ( .A0(n19349), .A1(y11[16]), .B0(n3026), .B1(temp2[16]), .Y(
        n19198) );
  OAI21XL U23441 ( .A0(n3063), .A1(n26554), .B0(n19198), .Y(n19435) );
  AOI22XL U23442 ( .A0(n19235), .A1(w2[49]), .B0(n19161), .B1(w1[81]), .Y(
        n19199) );
  INVX1 U23443 ( .A(n19438), .Y(n19901) );
  AOI22XL U23444 ( .A0(n19235), .A1(y11[17]), .B0(n19216), .B1(temp2[17]), .Y(
        n19200) );
  OAI21XL U23445 ( .A0(n3063), .A1(n26553), .B0(n19200), .Y(n19437) );
  AOI22XL U23446 ( .A0(n3027), .A1(w2[51]), .B0(n19161), .B1(w1[83]), .Y(
        n19202) );
  OAI21XL U23447 ( .A0(n19237), .A1(n25940), .B0(n19202), .Y(n19445) );
  AOI22XL U23448 ( .A0(n19235), .A1(y11[19]), .B0(n19216), .B1(temp2[19]), .Y(
        n19203) );
  OAI21XL U23449 ( .A0(n3063), .A1(n26551), .B0(n19203), .Y(n19444) );
  AOI22XL U23450 ( .A0(n19235), .A1(w2[50]), .B0(n19161), .B1(w1[82]), .Y(
        n19204) );
  OAI21XL U23451 ( .A0(n19237), .A1(n25890), .B0(n19204), .Y(n19442) );
  AOI22XL U23452 ( .A0(n19235), .A1(y11[18]), .B0(n19216), .B1(temp2[18]), .Y(
        n19205) );
  OAI21XL U23453 ( .A0(n3063), .A1(n26552), .B0(n19205), .Y(n19441) );
  NOR2XL U23454 ( .A(n19917), .B(n19441), .Y(n19206) );
  AOI22XL U23455 ( .A0(n3027), .A1(w2[52]), .B0(n19161), .B1(w1[84]), .Y(
        n19208) );
  OAI21XL U23456 ( .A0(n19237), .A1(n25939), .B0(n19208), .Y(n19426) );
  AOI22XL U23457 ( .A0(n19349), .A1(y11[20]), .B0(n19216), .B1(temp2[20]), .Y(
        n19209) );
  OAI21XL U23458 ( .A0(n3063), .A1(n26550), .B0(n19209), .Y(n19425) );
  NOR2XL U23459 ( .A(n19927), .B(n19425), .Y(n19212) );
  AOI22XL U23460 ( .A0(n3027), .A1(w2[53]), .B0(n19161), .B1(w1[85]), .Y(
        n19210) );
  OAI21XL U23461 ( .A0(n19237), .A1(n25889), .B0(n19210), .Y(n19428) );
  AOI22XL U23462 ( .A0(n19235), .A1(y11[21]), .B0(n19216), .B1(temp2[21]), .Y(
        n19211) );
  OAI21XL U23463 ( .A0(n3063), .A1(n26549), .B0(n19211), .Y(n19427) );
  AOI22XL U23464 ( .A0(n19346), .A1(w2[55]), .B0(n3026), .B1(w1[87]), .Y(
        n19213) );
  OAI21XL U23465 ( .A0(n19237), .A1(n26142), .B0(n19213), .Y(n19326) );
  AOI22XL U23466 ( .A0(n3027), .A1(w2[54]), .B0(n19161), .B1(w1[86]), .Y(
        n19215) );
  OAI21XL U23467 ( .A0(n19237), .A1(n25938), .B0(n19215), .Y(n19432) );
  AOI22XL U23468 ( .A0(n19235), .A1(y11[22]), .B0(n19216), .B1(temp2[22]), .Y(
        n19217) );
  OAI21XL U23469 ( .A0(n3063), .A1(n26548), .B0(n19217), .Y(n19431) );
  NOR2XL U23470 ( .A(n19937), .B(n19431), .Y(n19218) );
  AOI22XL U23471 ( .A0(n19349), .A1(w2[56]), .B0(n3062), .B1(w1[88]), .Y(
        n19221) );
  OAI21XL U23472 ( .A0(n3063), .A1(n26187), .B0(n19221), .Y(n19330) );
  AOI22XL U23473 ( .A0(y11[24]), .A1(n19346), .B0(n3062), .B1(temp2[24]), .Y(
        n19222) );
  OAI21XL U23474 ( .A0(n19237), .A1(n26510), .B0(n19222), .Y(n19329) );
  NOR2XL U23475 ( .A(n19265), .B(n19329), .Y(n19225) );
  OAI21XL U23476 ( .A0(n3063), .A1(n25936), .B0(n19223), .Y(n19334) );
  AOI22XL U23477 ( .A0(y11[25]), .A1(n19235), .B0(n3062), .B1(temp2[25]), .Y(
        n19224) );
  OAI21XL U23478 ( .A0(n3063), .A1(n26511), .B0(n19224), .Y(n19333) );
  NOR2XL U23479 ( .A(n19301), .B(n19333), .Y(n19268) );
  AOI22XL U23480 ( .A0(n3027), .A1(w2[59]), .B0(n3062), .B1(w1[91]), .Y(n19226) );
  OAI21XL U23481 ( .A0(n3063), .A1(n25937), .B0(n19226), .Y(n19311) );
  AOI22XL U23482 ( .A0(y11[27]), .A1(n19235), .B0(n19216), .B1(temp2[27]), .Y(
        n19227) );
  OAI21XL U23483 ( .A0(n3063), .A1(n26512), .B0(n19227), .Y(n19310) );
  AOI22XL U23484 ( .A0(n19349), .A1(w2[58]), .B0(n19161), .B1(w1[90]), .Y(
        n19228) );
  OAI21XL U23485 ( .A0(n19237), .A1(n26185), .B0(n19228), .Y(n19338) );
  OAI21XL U23486 ( .A0(n19237), .A1(n26505), .B0(n19229), .Y(n19337) );
  AOI22XL U23487 ( .A0(n3027), .A1(w2[60]), .B0(n3062), .B1(w1[92]), .Y(n19232) );
  OAI21XL U23488 ( .A0(n19237), .A1(n26186), .B0(n19232), .Y(n19315) );
  AOI22XL U23489 ( .A0(y11[28]), .A1(n19235), .B0(n19216), .B1(temp2[28]), .Y(
        n19233) );
  OAI21XL U23490 ( .A0(n19237), .A1(n26506), .B0(n19233), .Y(n19314) );
  NOR2XL U23491 ( .A(n19294), .B(n19314), .Y(n19238) );
  AOI22XL U23492 ( .A0(n19349), .A1(w2[61]), .B0(n3062), .B1(w1[93]), .Y(
        n19234) );
  OAI21XL U23493 ( .A0(n19237), .A1(n25935), .B0(n19234), .Y(n19319) );
  AOI22XL U23494 ( .A0(y11[29]), .A1(n19235), .B0(n3062), .B1(temp2[29]), .Y(
        n19236) );
  OAI21XL U23495 ( .A0(n19237), .A1(n26508), .B0(n19236), .Y(n19318) );
  NAND2XL U23496 ( .A(n19841), .B(n19435), .Y(n19244) );
  NAND2XL U23497 ( .A(n19901), .B(n19437), .Y(n19243) );
  OAI21XL U23498 ( .A0(n19245), .A1(n19244), .B0(n19243), .Y(n19250) );
  NAND2XL U23499 ( .A(n19917), .B(n19441), .Y(n19247) );
  NAND2XL U23500 ( .A(n19922), .B(n19444), .Y(n19246) );
  OAI21XL U23501 ( .A0(n19248), .A1(n19247), .B0(n19246), .Y(n19249) );
  AOI21XL U23502 ( .A0(n19251), .A1(n19250), .B0(n19249), .Y(n19264) );
  NAND2XL U23503 ( .A(n19927), .B(n19425), .Y(n19253) );
  NAND2XL U23504 ( .A(n19932), .B(n19427), .Y(n19252) );
  OAI21XL U23505 ( .A0(n19254), .A1(n19253), .B0(n19252), .Y(n19260) );
  NAND2XL U23506 ( .A(n19937), .B(n19431), .Y(n19257) );
  NAND2XL U23507 ( .A(n19255), .B(n19325), .Y(n19256) );
  OAI21XL U23508 ( .A0(n19258), .A1(n19257), .B0(n19256), .Y(n19259) );
  AOI21XL U23509 ( .A0(n19261), .A1(n19260), .B0(n19259), .Y(n19262) );
  NAND2XL U23510 ( .A(n19265), .B(n19329), .Y(n19267) );
  NAND2XL U23511 ( .A(n19301), .B(n19333), .Y(n19266) );
  OAI21XL U23512 ( .A0(n19268), .A1(n19267), .B0(n19266), .Y(n19273) );
  NAND2XL U23513 ( .A(n19299), .B(n19337), .Y(n19270) );
  NAND2XL U23514 ( .A(n19296), .B(n19310), .Y(n19269) );
  OAI21XL U23515 ( .A0(n19271), .A1(n19270), .B0(n19269), .Y(n19272) );
  AOI21XL U23516 ( .A0(n19274), .A1(n19273), .B0(n19272), .Y(n19283) );
  NAND2XL U23517 ( .A(n19294), .B(n19314), .Y(n19276) );
  NAND2XL U23518 ( .A(n19292), .B(n19318), .Y(n19275) );
  OAI21XL U23519 ( .A0(n19277), .A1(n19276), .B0(n19275), .Y(n19280) );
  INVX4 U23520 ( .A(n19297), .Y(n19564) );
  OAI21X2 U23521 ( .A0(n19566), .A1(n19292), .B0(n19291), .Y(n24433) );
  NAND2XL U23522 ( .A(n19564), .B(n19310), .Y(n19295) );
  OAI21X2 U23523 ( .A0(n19566), .A1(n19265), .B0(n19302), .Y(n24092) );
  OAI21X2 U23524 ( .A0(n19566), .A1(n19255), .B0(n19303), .Y(n24309) );
  CMPR22X1 U23525 ( .A(n24433), .B(n19304), .CO(n20130), .S(n24435) );
  CMPR22X1 U23526 ( .A(n24390), .B(n19305), .CO(n19304), .S(n24391) );
  CMPR22X1 U23527 ( .A(n24295), .B(n19306), .CO(n19305), .S(n24296) );
  NAND2XL U23528 ( .A(n19564), .B(n19311), .Y(n19312) );
  OAI21XL U23529 ( .A0(n19564), .A1(n19313), .B0(n19312), .Y(n23206) );
  OAI21XL U23530 ( .A0(n19564), .A1(n19107), .B0(n19324), .Y(n23203) );
  NAND2XL U23531 ( .A(n3041), .B(n19326), .Y(n19327) );
  NAND2XL U23532 ( .A(n3041), .B(n19338), .Y(n19339) );
  NOR2X1 U23533 ( .A(n24309), .B(n19363), .Y(n19361) );
  INVXL U23534 ( .A(n19399), .Y(n19355) );
  INVXL U23535 ( .A(n19358), .Y(n19360) );
  NAND2XL U23536 ( .A(n19360), .B(n19359), .Y(n19362) );
  XOR2X1 U23537 ( .A(n19362), .B(n19361), .Y(n19457) );
  XNOR2X1 U23538 ( .A(n24309), .B(n19363), .Y(n19510) );
  NAND2XL U23539 ( .A(n3039), .B(n19368), .Y(n19369) );
  OAI21XL U23540 ( .A0(n3039), .A1(n19659), .B0(n19369), .Y(n19481) );
  OAI21XL U23541 ( .A0(n19564), .A1(n19816), .B0(n19372), .Y(n19663) );
  OAI21XL U23542 ( .A0(n19564), .A1(n19821), .B0(n19375), .Y(n19649) );
  NAND2XL U23543 ( .A(n3039), .B(n19649), .Y(n19376) );
  OAI21XL U23544 ( .A0(n3039), .A1(n19377), .B0(n19376), .Y(n19500) );
  INVXL U23545 ( .A(n19500), .Y(n19378) );
  NAND2XL U23546 ( .A(n3035), .B(n19378), .Y(n19379) );
  OAI21XL U23547 ( .A0(n19457), .A1(n19481), .B0(n19379), .Y(n19740) );
  INVXL U23548 ( .A(n19396), .Y(n19380) );
  NAND2XL U23549 ( .A(n19380), .B(n19398), .Y(n19381) );
  OAI21XL U23550 ( .A0(n19566), .A1(n19480), .B0(n19387), .Y(n19669) );
  NAND2XL U23551 ( .A(n3039), .B(n19669), .Y(n19388) );
  OAI21XL U23552 ( .A0(n3039), .A1(n19627), .B0(n19388), .Y(n19489) );
  OAI21XL U23553 ( .A0(n19564), .A1(n19788), .B0(n19391), .Y(n19622) );
  OAI21XL U23554 ( .A0(n19564), .A1(n19795), .B0(n19394), .Y(n19648) );
  AOI22XL U23555 ( .A0(n3094), .A1(n19622), .B0(n3039), .B1(n19648), .Y(n19483) );
  NAND2XL U23556 ( .A(n3035), .B(n19483), .Y(n19395) );
  OAI21XL U23557 ( .A0(n19457), .A1(n19489), .B0(n19395), .Y(n19743) );
  OAI22XL U23558 ( .A0(n19740), .A1(n3036), .B0(n19542), .B1(n19743), .Y(
        n19576) );
  NOR2XL U23559 ( .A(n19396), .B(n19399), .Y(n19402) );
  OAI21XL U23560 ( .A0(n19399), .A1(n19398), .B0(n19397), .Y(n19400) );
  OAI21XL U23561 ( .A0(n19423), .A1(n19419), .B0(n19420), .Y(n19408) );
  NAND2XL U23562 ( .A(n24390), .B(n19404), .Y(n19405) );
  INVXL U23563 ( .A(n19419), .Y(n19421) );
  NAND2XL U23564 ( .A(n3039), .B(n19643), .Y(n19430) );
  OAI21XL U23565 ( .A0(n3039), .A1(n19623), .B0(n19430), .Y(n19493) );
  OAI21XL U23566 ( .A0(n3041), .A1(n19938), .B0(n19433), .Y(n19642) );
  NAND2XL U23567 ( .A(n3035), .B(n19502), .Y(n19434) );
  OAI21XL U23568 ( .A0(n3035), .A1(n19493), .B0(n19434), .Y(n19797) );
  INVXL U23569 ( .A(n19797), .Y(n19451) );
  OAI21XL U23570 ( .A0(n19564), .A1(n19902), .B0(n19439), .Y(n19615) );
  NAND2XL U23571 ( .A(n3039), .B(n19615), .Y(n19440) );
  OAI21XL U23572 ( .A0(n3039), .A1(n19676), .B0(n19440), .Y(n19497) );
  OAI21XL U23573 ( .A0(n19564), .A1(n19918), .B0(n19443), .Y(n19641) );
  NAND2XL U23574 ( .A(n3039), .B(n19625), .Y(n19447) );
  OAI21XL U23575 ( .A0(n3039), .A1(n19448), .B0(n19447), .Y(n19496) );
  INVXL U23576 ( .A(n19496), .Y(n19449) );
  NAND2XL U23577 ( .A(n3035), .B(n19449), .Y(n19450) );
  OAI21XL U23578 ( .A0(n3035), .A1(n19497), .B0(n19450), .Y(n19741) );
  AOI22XL U23579 ( .A0(n3094), .A1(n19669), .B0(n3039), .B1(n19622), .Y(n19525) );
  NAND2XL U23580 ( .A(n3039), .B(n19458), .Y(n19459) );
  OAI21XL U23581 ( .A0(n3039), .A1(n19460), .B0(n19459), .Y(n19521) );
  INVXL U23582 ( .A(n19521), .Y(n19461) );
  AOI22XL U23583 ( .A0(n3166), .A1(n19525), .B0(n19461), .B1(n3035), .Y(n19543) );
  NAND2XL U23584 ( .A(n3039), .B(n19663), .Y(n19462) );
  OAI21XL U23585 ( .A0(n3039), .A1(n19646), .B0(n19462), .Y(n19518) );
  AOI22XL U23586 ( .A0(n3094), .A1(n19649), .B0(n3039), .B1(n19463), .Y(n19513) );
  NAND2XL U23587 ( .A(n3035), .B(n19513), .Y(n19464) );
  OAI21XL U23588 ( .A0(n3035), .A1(n19518), .B0(n19464), .Y(n19535) );
  NAND2XL U23589 ( .A(n3039), .B(n19642), .Y(n19465) );
  OAI21XL U23590 ( .A0(n3039), .A1(n19466), .B0(n19465), .Y(n19514) );
  OAI21XL U23591 ( .A0(n3035), .A1(n19514), .B0(n19467), .Y(n19804) );
  INVXL U23592 ( .A(n19804), .Y(n19475) );
  NAND2XL U23593 ( .A(n3039), .B(n19641), .Y(n19468) );
  OAI21XL U23594 ( .A0(n3039), .A1(n19469), .B0(n19468), .Y(n19511) );
  NAND2XL U23595 ( .A(n3039), .B(n19470), .Y(n19471) );
  OAI21XL U23596 ( .A0(n3039), .A1(n19472), .B0(n19471), .Y(n19517) );
  INVXL U23597 ( .A(n19517), .Y(n19473) );
  NAND2XL U23598 ( .A(n3035), .B(n19473), .Y(n19474) );
  OAI21XL U23599 ( .A0(n3035), .A1(n19511), .B0(n19474), .Y(n19536) );
  OAI21XL U23600 ( .A0(n3165), .A1(n19478), .B0(n19477), .Y(n19777) );
  INVXL U23601 ( .A(n19481), .Y(n19482) );
  AOI22XL U23602 ( .A0(n3166), .A1(n19483), .B0(n19482), .B1(n3035), .Y(n19712) );
  NAND2XL U23603 ( .A(n19564), .B(n19487), .Y(n19488) );
  OAI21XL U23604 ( .A0(n19566), .A1(n19533), .B0(n19488), .Y(n19630) );
  AOI22XL U23605 ( .A0(n3094), .A1(n19666), .B0(n3039), .B1(n19630), .Y(n19570) );
  INVXL U23606 ( .A(n19570), .Y(n19492) );
  INVXL U23607 ( .A(n19489), .Y(n19490) );
  NAND2XL U23608 ( .A(n3035), .B(n19490), .Y(n19491) );
  OAI21XL U23609 ( .A0(n3035), .A1(n19492), .B0(n19491), .Y(n19708) );
  AOI2BB2XL U23610 ( .B0(n19712), .B1(n19542), .A0N(n19542), .A1N(n19708), .Y(
        n19608) );
  INVXL U23611 ( .A(n19493), .Y(n19494) );
  NAND2XL U23612 ( .A(n3035), .B(n19494), .Y(n19495) );
  OAI21XL U23613 ( .A0(n3035), .A1(n19496), .B0(n19495), .Y(n19713) );
  INVXL U23614 ( .A(n19713), .Y(n19501) );
  INVXL U23615 ( .A(n19497), .Y(n19498) );
  NAND2XL U23616 ( .A(n3035), .B(n19498), .Y(n19499) );
  OAI21XL U23617 ( .A0(n3035), .A1(n19500), .B0(n19499), .Y(n19711) );
  AOI22XL U23618 ( .A0(n19504), .A1(n19503), .B0(n19730), .B1(n19934), .Y(
        n19505) );
  NAND2XL U23619 ( .A(n4622), .B(n3166), .Y(n19644) );
  INVXL U23620 ( .A(n19511), .Y(n19512) );
  AOI22XL U23621 ( .A0(n3166), .A1(n19513), .B0(n19512), .B1(n3035), .Y(n19727) );
  INVXL U23622 ( .A(n19514), .Y(n19515) );
  NAND2XL U23623 ( .A(n3035), .B(n19515), .Y(n19516) );
  OAI21XL U23624 ( .A0(n3035), .A1(n19517), .B0(n19516), .Y(n19728) );
  INVXL U23625 ( .A(n19518), .Y(n19519) );
  NAND2XL U23626 ( .A(n3035), .B(n19519), .Y(n19520) );
  OAI21XL U23627 ( .A0(n3035), .A1(n19521), .B0(n19520), .Y(n19726) );
  INVXL U23628 ( .A(n19630), .Y(n19524) );
  NAND2XL U23629 ( .A(n3039), .B(n19522), .Y(n19523) );
  OAI21XL U23630 ( .A0(n3039), .A1(n19524), .B0(n19523), .Y(n19540) );
  NAND2XL U23631 ( .A(n3035), .B(n19525), .Y(n19526) );
  OAI21XL U23632 ( .A0(n3035), .A1(n19540), .B0(n19526), .Y(n19722) );
  OAI22XL U23633 ( .A0(n19726), .A1(n3036), .B0(n19542), .B1(n19722), .Y(
        n19696) );
  OAI21XL U23634 ( .A0(n19696), .A1(n19807), .B0(n19747), .Y(n19527) );
  INVXL U23635 ( .A(n19748), .Y(n19580) );
  NAND2X1 U23636 ( .A(n2996), .B(n4622), .Y(n19739) );
  NAND2XL U23637 ( .A(n19564), .B(n19538), .Y(n19539) );
  OAI21XL U23638 ( .A0(n19566), .A1(n19552), .B0(n19539), .Y(n19652) );
  AOI22XL U23639 ( .A0(n3094), .A1(n19652), .B0(n3039), .B1(n19666), .Y(n19689) );
  INVXL U23640 ( .A(n19540), .Y(n19541) );
  AOI22XL U23641 ( .A0(n3166), .A1(n19689), .B0(n19541), .B1(n3035), .Y(n19588) );
  OAI21XL U23642 ( .A0(n19806), .A1(n2996), .B0(n19545), .Y(n19546) );
  INVXL U23643 ( .A(n19838), .Y(n19578) );
  INVXL U23644 ( .A(n19665), .Y(n19559) );
  INVXL U23645 ( .A(n19661), .Y(n19558) );
  AOI22XL U23646 ( .A0(n3094), .A1(n19559), .B0(n3039), .B1(n19558), .Y(n19602) );
  NAND2XL U23647 ( .A(n19564), .B(n19563), .Y(n19565) );
  OAI21XL U23648 ( .A0(n19564), .A1(n19737), .B0(n19565), .Y(n19634) );
  AOI22XL U23649 ( .A0(n3094), .A1(n19650), .B0(n3039), .B1(n19634), .Y(n19605) );
  AOI22XL U23650 ( .A0(n3166), .A1(n19602), .B0(n19605), .B1(n3035), .Y(n19573) );
  NAND2XL U23651 ( .A(n3039), .B(n19652), .Y(n19569) );
  OAI21XL U23652 ( .A0(n3039), .A1(n19632), .B0(n19569), .Y(n19603) );
  NAND2XL U23653 ( .A(n3035), .B(n19570), .Y(n19571) );
  OAI21XL U23654 ( .A0(n3035), .A1(n19603), .B0(n19571), .Y(n19742) );
  INVXL U23655 ( .A(n19742), .Y(n19572) );
  AOI22XL U23656 ( .A0(n19573), .A1(n3036), .B0(n19572), .B1(n19542), .Y(
        n19574) );
  AOI21XL U23657 ( .A0(n19574), .A1(n3159), .B0(n19730), .Y(n19575) );
  OAI21XL U23658 ( .A0(n2996), .A1(n19576), .B0(n19575), .Y(n19577) );
  OAI21XL U23659 ( .A0(n19578), .A1(n19747), .B0(n19577), .Y(n19579) );
  NAND2XL U23660 ( .A(n19580), .B(n19579), .Y(n19582) );
  AOI21XL U23661 ( .A0(n19582), .A1(n19952), .B0(n3164), .Y(n19581) );
  OAI21XL U23662 ( .A0(n3165), .A1(n19582), .B0(n19581), .Y(n19702) );
  NAND2XL U23663 ( .A(n3039), .B(n19650), .Y(n19585) );
  OAI21XL U23664 ( .A0(n3039), .A1(n19661), .B0(n19585), .Y(n19691) );
  INVXL U23665 ( .A(n19691), .Y(n19587) );
  INVXL U23666 ( .A(n19632), .Y(n19586) );
  AOI22XL U23667 ( .A0(n3094), .A1(n19634), .B0(n3039), .B1(n19586), .Y(n19690) );
  AOI22XL U23668 ( .A0(n3166), .A1(n19587), .B0(n19690), .B1(n3035), .Y(n19589) );
  AOI22XL U23669 ( .A0(n19589), .A1(n3036), .B0(n19588), .B1(n19542), .Y(
        n19590) );
  AOI21XL U23670 ( .A0(n19590), .A1(n3159), .B0(n19730), .Y(n19594) );
  NAND2XL U23671 ( .A(n19591), .B(n19807), .Y(n19593) );
  AOI22XL U23672 ( .A0(n19594), .A1(n19593), .B0(n19898), .B1(n19730), .Y(
        n19595) );
  AOI21XL U23673 ( .A0(n19597), .A1(n19952), .B0(n3164), .Y(n19596) );
  OAI21XL U23674 ( .A0(n3165), .A1(n19597), .B0(n19596), .Y(n19704) );
  OR2X2 U23675 ( .A(n19704), .B(n19703), .Y(n20037) );
  NAND2XL U23676 ( .A(n20069), .B(n20037), .Y(n19707) );
  AOI22XL U23677 ( .A0(n19601), .A1(n3159), .B0(n19807), .B1(n19600), .Y(
        n19812) );
  NOR2XL U23678 ( .A(n3166), .B(n19602), .Y(n19606) );
  INVXL U23679 ( .A(n19603), .Y(n19604) );
  AOI22XL U23680 ( .A0(n3166), .A1(n19605), .B0(n19604), .B1(n3035), .Y(n19709) );
  AOI22XL U23681 ( .A0(n19606), .A1(n3036), .B0(n19709), .B1(n19542), .Y(
        n19607) );
  AOI21XL U23682 ( .A0(n19607), .A1(n3159), .B0(n19730), .Y(n19610) );
  NAND2XL U23683 ( .A(n19608), .B(n19807), .Y(n19609) );
  AOI22XL U23684 ( .A0(n19730), .A1(n19812), .B0(n19610), .B1(n19609), .Y(
        n19611) );
  NOR2XL U23685 ( .A(n19611), .B(n19748), .Y(n19613) );
  NAND2XL U23686 ( .A(n19613), .B(n19796), .Y(n19612) );
  OAI211XL U23687 ( .A0(n3215), .A1(n19613), .B0(n6192), .C0(n19612), .Y(
        n19614) );
  NAND2XL U23688 ( .A(n3166), .B(n3094), .Y(n19664) );
  NAND2XL U23689 ( .A(n19542), .B(n19664), .Y(n19640) );
  OAI21XL U23690 ( .A0(n2996), .A1(n19640), .B0(n19747), .Y(n19621) );
  NAND2XL U23691 ( .A(n19739), .B(n19615), .Y(n19618) );
  AOI31XL U23692 ( .A0(n19618), .A1(n19617), .A2(n19616), .B0(n19747), .Y(
        n19620) );
  AOI211XL U23693 ( .A0(n19622), .A1(n19621), .B0(n19620), .C0(n19619), .Y(
        n19639) );
  INVXL U23694 ( .A(n19739), .Y(n19678) );
  AOI211XL U23695 ( .A0(n3159), .A1(n3166), .B0(n19678), .C0(n19747), .Y(
        n19624) );
  OAI21XL U23696 ( .A0(n19626), .A1(n19625), .B0(n19624), .Y(n19638) );
  NOR2XL U23697 ( .A(n19730), .B(n19542), .Y(n19628) );
  AOI21XL U23698 ( .A0(n19628), .A1(n3094), .B0(n19627), .Y(n19631) );
  AOI21XL U23699 ( .A0(n19628), .A1(n3166), .B0(n19662), .Y(n19629) );
  OAI21XL U23700 ( .A0(n19631), .A1(n19630), .B0(n19629), .Y(n19637) );
  AOI21XL U23701 ( .A0(n19662), .A1(n3094), .B0(n19632), .Y(n19635) );
  OAI21XL U23702 ( .A0(n3036), .A1(n3166), .B0(n19662), .Y(n19633) );
  OAI21XL U23703 ( .A0(n19635), .A1(n19634), .B0(n19633), .Y(n19636) );
  NAND4XL U23704 ( .A(n19639), .B(n19638), .C(n19637), .D(n19636), .Y(n19685)
         );
  INVXL U23705 ( .A(n19664), .Y(n19729) );
  OAI21XL U23706 ( .A0(n19644), .A1(n19643), .B0(n19807), .Y(n19645) );
  AOI31XL U23707 ( .A0(n19647), .A1(n19646), .A2(n19645), .B0(n19747), .Y(
        n19657) );
  AOI21XL U23708 ( .A0(n19678), .A1(n3166), .B0(n19747), .Y(n19675) );
  NAND2XL U23709 ( .A(n19807), .B(n19542), .Y(n19668) );
  OAI21XL U23710 ( .A0(n19668), .A1(n3166), .B0(n19747), .Y(n19658) );
  AOI22XL U23711 ( .A0(n19675), .A1(n19649), .B0(n19658), .B1(n19648), .Y(
        n19656) );
  INVXL U23712 ( .A(n19662), .Y(n19653) );
  AOI22XL U23713 ( .A0(n19653), .A1(n19652), .B0(n19651), .B1(n19650), .Y(
        n19655) );
  NAND4BXL U23714 ( .AN(n19657), .B(n19656), .C(n19655), .D(n19654), .Y(n19682) );
  INVXL U23715 ( .A(n19658), .Y(n19660) );
  AOI211XL U23716 ( .A0(n19747), .A1(n3094), .B0(n19660), .C0(n19659), .Y(
        n19681) );
  AOI22XL U23717 ( .A0(n19662), .A1(n3036), .B0(n19661), .B1(n19665), .Y(
        n19674) );
  OAI211XL U23718 ( .A0(n19664), .A1(n19739), .B0(n19730), .C0(n19663), .Y(
        n19673) );
  AOI22XL U23719 ( .A0(n19667), .A1(n19666), .B0(n19692), .B1(n3035), .Y(
        n19672) );
  INVXL U23720 ( .A(n19668), .Y(n19670) );
  OAI21XL U23721 ( .A0(n19670), .A1(n19730), .B0(n19669), .Y(n19671) );
  INVXL U23722 ( .A(n19675), .Y(n19677) );
  AOI211XL U23723 ( .A0(n19678), .A1(n3094), .B0(n19677), .C0(n19676), .Y(
        n19679) );
  OR4X2 U23724 ( .A(n19682), .B(n19679), .C(n19680), .D(n19681), .Y(n19684) );
  AOI22XL U23725 ( .A0(n19688), .A1(n19807), .B0(n19687), .B1(n3159), .Y(
        n19817) );
  NAND2XL U23726 ( .A(n19817), .B(n19730), .Y(n19698) );
  AOI22XL U23727 ( .A0(n3166), .A1(n19690), .B0(n19689), .B1(n3035), .Y(n19724) );
  AOI22XL U23728 ( .A0(n3166), .A1(n19692), .B0(n19457), .B1(n19691), .Y(
        n19693) );
  AOI21XL U23729 ( .A0(n19694), .A1(n3159), .B0(n19730), .Y(n19695) );
  OAI21XL U23730 ( .A0(n2996), .A1(n19696), .B0(n19695), .Y(n19697) );
  AOI21XL U23731 ( .A0(n19698), .A1(n19697), .B0(n19748), .Y(n19700) );
  NAND2XL U23732 ( .A(n19700), .B(n19796), .Y(n19699) );
  OAI211XL U23733 ( .A0(n19700), .A1(n3215), .B0(n6192), .C0(n19699), .Y(
        n20072) );
  NAND2XL U23734 ( .A(n19702), .B(n19701), .Y(n20068) );
  INVXL U23735 ( .A(n20068), .Y(n20035) );
  NAND2XL U23736 ( .A(n19704), .B(n19703), .Y(n20036) );
  INVXL U23737 ( .A(n20036), .Y(n19705) );
  AOI21XL U23738 ( .A0(n20037), .A1(n20035), .B0(n19705), .Y(n19706) );
  AOI21XL U23739 ( .A0(n19710), .A1(n3159), .B0(n19730), .Y(n19716) );
  NAND2XL U23740 ( .A(n19783), .B(n19807), .Y(n19715) );
  OAI21XL U23741 ( .A0(n3165), .A1(n19719), .B0(n19718), .Y(n19755) );
  NOR2XL U23742 ( .A(n19755), .B(n19754), .Y(n20026) );
  INVXL U23743 ( .A(n20026), .Y(n20031) );
  INVXL U23744 ( .A(n19722), .Y(n19723) );
  AOI22XL U23745 ( .A0(n19724), .A1(n3036), .B0(n19723), .B1(n19542), .Y(
        n19725) );
  AOI21XL U23746 ( .A0(n19725), .A1(n3159), .B0(n19730), .Y(n19732) );
  NAND2XL U23747 ( .A(n19790), .B(n19807), .Y(n19731) );
  AOI22XL U23748 ( .A0(n19732), .A1(n19731), .B0(n19919), .B1(n19730), .Y(
        n19733) );
  AOI21XL U23749 ( .A0(n19735), .A1(n19952), .B0(n3164), .Y(n19734) );
  OAI21XL U23750 ( .A0(n3165), .A1(n19735), .B0(n19734), .Y(n19757) );
  NAND2XL U23751 ( .A(n20031), .B(n19738), .Y(n20020) );
  OAI22XL U23752 ( .A0(n19741), .A1(n3036), .B0(n19542), .B1(n19740), .Y(
        n19799) );
  OAI22XL U23753 ( .A0(n19743), .A1(n3036), .B0(n19542), .B1(n19742), .Y(
        n19744) );
  OAI22XL U23754 ( .A0(n19799), .A1(n2996), .B0(n19744), .B1(n19807), .Y(
        n19745) );
  NAND2XL U23755 ( .A(n19745), .B(n19747), .Y(n19746) );
  OAI21XL U23756 ( .A0(n19924), .A1(n19747), .B0(n19746), .Y(n19749) );
  AOI21XL U23757 ( .A0(n19751), .A1(n19952), .B0(n3164), .Y(n19750) );
  OAI21XL U23758 ( .A0(n3165), .A1(n19751), .B0(n19750), .Y(n19761) );
  NOR2XL U23759 ( .A(n19761), .B(n19760), .Y(n20021) );
  NOR2XL U23760 ( .A(n20020), .B(n20021), .Y(n19763) );
  NAND2XL U23761 ( .A(n19755), .B(n19754), .Y(n20030) );
  INVXL U23762 ( .A(n20030), .Y(n19759) );
  NAND2XL U23763 ( .A(n19757), .B(n19756), .Y(n20027) );
  INVXL U23764 ( .A(n20027), .Y(n19758) );
  NAND2XL U23765 ( .A(n19761), .B(n19760), .Y(n20022) );
  OAI21XL U23766 ( .A0(n20019), .A1(n20021), .B0(n20022), .Y(n19762) );
  OAI21XL U23767 ( .A0(n19773), .A1(n20055), .B0(n19772), .Y(n20046) );
  OAI21XL U23768 ( .A0(n19892), .A1(n20049), .B0(n19893), .Y(n19778) );
  OAI21XL U23769 ( .A0(n19542), .A1(n19797), .B0(n19807), .Y(n19798) );
  OAI21XL U23770 ( .A0(n3165), .A1(n19801), .B0(n19800), .Y(n19827) );
  OAI21XL U23771 ( .A0(n19542), .A1(n19804), .B0(n19807), .Y(n19805) );
  OAI21XL U23772 ( .A0(n3165), .A1(n19809), .B0(n19808), .Y(n19829) );
  OAI21XL U23773 ( .A0(n3165), .A1(n19814), .B0(n19813), .Y(n19833) );
  OAI21XL U23774 ( .A0(n3165), .A1(n19819), .B0(n19818), .Y(n19835) );
  OAI21XL U23775 ( .A0(n19878), .A1(n19884), .B0(n19879), .Y(n19871) );
  OAI21XL U23776 ( .A0(n19865), .A1(n19874), .B0(n19866), .Y(n19830) );
  OAI21XL U23777 ( .A0(n19852), .A1(n19857), .B0(n19853), .Y(n19983) );
  AOI21XL U23778 ( .A0(n19989), .A1(n19980), .B0(n19983), .Y(n19836) );
  OAI21XL U23779 ( .A0(n19992), .A1(n19837), .B0(n19836), .Y(n19847) );
  OAI21XL U23780 ( .A0(n3165), .A1(n19840), .B0(n19839), .Y(n19844) );
  OAI21XL U23781 ( .A0(n19992), .A1(n19851), .B0(n19850), .Y(n19856) );
  OAI21XL U23782 ( .A0(n19992), .A1(n19903), .B0(n19910), .Y(n19860) );
  AOI21XL U23783 ( .A0(n19871), .A1(n19875), .B0(n19862), .Y(n19863) );
  OAI21XL U23784 ( .A0(n19992), .A1(n19864), .B0(n19863), .Y(n19869) );
  OAI21XL U23785 ( .A0(n19992), .A1(n19873), .B0(n19872), .Y(n19877) );
  XNOR2X1 U23786 ( .A(n19877), .B(n19876), .Y(n20254) );
  OAI21XL U23787 ( .A0(n19992), .A1(n19883), .B0(n19884), .Y(n19882) );
  NOR2X1 U23788 ( .A(n20254), .B(n20255), .Y(n20110) );
  XOR2X1 U23789 ( .A(n19992), .B(n19886), .Y(n20235) );
  OAI21XL U23790 ( .A0(n19889), .A1(n20048), .B0(n20049), .Y(n19890) );
  OAI21XL U23791 ( .A0(n3165), .A1(n19900), .B0(n19899), .Y(n19905) );
  OAI21XL U23792 ( .A0(n19993), .A1(n19984), .B0(n19994), .Y(n19906) );
  OAI21XL U23793 ( .A0(n3165), .A1(n19916), .B0(n19915), .Y(n19940) );
  OAI21XL U23794 ( .A0(n3165), .A1(n19921), .B0(n19920), .Y(n19942) );
  OR2X2 U23795 ( .A(n19999), .B(n19959), .Y(n19963) );
  OAI21XL U23796 ( .A0(n20012), .A1(n20005), .B0(n20013), .Y(n19947) );
  OAI21XL U23797 ( .A0(n19998), .A1(n19959), .B0(n19955), .Y(n19956) );
  OAI21XL U23798 ( .A0(n20011), .A1(n19967), .B0(n19966), .Y(n19970) );
  OAI21XL U23799 ( .A0(n20011), .A1(n19976), .B0(n19977), .Y(n19975) );
  OAI21XL U23800 ( .A0(n19986), .A1(n19985), .B0(n19984), .Y(n19987) );
  OAI21XL U23801 ( .A0(n19992), .A1(n19991), .B0(n19990), .Y(n19997) );
  OAI21XL U23802 ( .A0(n20011), .A1(n19999), .B0(n19998), .Y(n20003) );
  AOI21XL U23803 ( .A0(n20008), .A1(n20007), .B0(n20006), .Y(n20009) );
  OAI21XL U23804 ( .A0(n20011), .A1(n20010), .B0(n20009), .Y(n20016) );
  CMPR22X1 U23805 ( .A(n24072), .B(n20017), .CO(n19306), .S(n24073) );
  OAI21XL U23806 ( .A0(n20033), .A1(n20020), .B0(n20019), .Y(n20025) );
  OAI21XL U23807 ( .A0(n20033), .A1(n20026), .B0(n20030), .Y(n20029) );
  NAND2XL U23808 ( .A(n19738), .B(n20027), .Y(n20028) );
  XNOR2X1 U23809 ( .A(n20029), .B(n20028), .Y(n20199) );
  NAND2XL U23810 ( .A(n20031), .B(n20030), .Y(n20032) );
  XOR2X1 U23811 ( .A(n20033), .B(n20032), .Y(n20203) );
  INVXL U23812 ( .A(n20034), .Y(n20071) );
  NAND2XL U23813 ( .A(n20037), .B(n20036), .Y(n20038) );
  XOR2X1 U23814 ( .A(n20039), .B(n20038), .Y(n20204) );
  AOI21XL U23815 ( .A0(n20059), .A1(n20044), .B0(n20040), .Y(n20043) );
  AOI21XL U23816 ( .A0(n20059), .A1(n20047), .B0(n20046), .Y(n20052) );
  OAI21XL U23817 ( .A0(n20056), .A1(n20055), .B0(n20054), .Y(n20057) );
  AOI21XL U23818 ( .A0(n20059), .A1(n20058), .B0(n20057), .Y(n20062) );
  OR2X2 U23819 ( .A(n20188), .B(n20186), .Y(n20107) );
  CMPR22X1 U23820 ( .A(n24341), .B(n20067), .CO(n20017), .S(n24342) );
  NAND2XL U23821 ( .A(n20069), .B(n20068), .Y(n20070) );
  INVXL U23822 ( .A(n20072), .Y(n20073) );
  OAI21XL U23823 ( .A0(n20077), .A1(n20076), .B0(n20075), .Y(n20079) );
  AOI31X1 U23824 ( .A0(n20111), .A1(n20082), .A2(n20114), .B0(n20081), .Y(
        n24894) );
  AOI2BB1XL U23825 ( .A0N(n20084), .A1N(n20199), .B0(n20177), .Y(n20085) );
  AOI2BB1XL U23826 ( .A0N(n20196), .A1N(n20085), .B0(n20195), .Y(n20086) );
  AOI2BB1XL U23827 ( .A0N(n20086), .A1N(n20186), .B0(n20188), .Y(n20087) );
  INVXL U23828 ( .A(n20236), .Y(n20088) );
  AOI2BB1XL U23829 ( .A0N(n20090), .A1N(n20255), .B0(n20254), .Y(n20091) );
  INVXL U23830 ( .A(n24680), .Y(n20092) );
  AOI2BB1X1 U23831 ( .A0N(n20094), .A1N(n24716), .B0(n24798), .Y(n20095) );
  INVXL U23832 ( .A(n24828), .Y(n20096) );
  AOI2BB1X2 U23833 ( .A0N(n20098), .A1N(n24889), .B0(n24938), .Y(n20099) );
  INVXL U23834 ( .A(n24937), .Y(n20100) );
  AOI21X1 U23835 ( .A0(n20101), .A1(n20100), .B0(n25344), .Y(n20102) );
  AOI2BB1X2 U23836 ( .A0N(n20102), .A1N(n25343), .B0(n20167), .Y(n20125) );
  OAI21XL U23837 ( .A0(n20156), .A1(n24063), .B0(n20103), .Y(n20104) );
  OAI21XL U23838 ( .A0(n20108), .A1(n20107), .B0(n20106), .Y(n20109) );
  CMPR22X1 U23839 ( .A(n24092), .B(n24309), .CO(n20067), .S(n24093) );
  XOR2X1 U23840 ( .A(n24435), .B(n20119), .Y(n24432) );
  INVXL U23841 ( .A(n24391), .Y(n20120) );
  CMPR32X1 U23842 ( .A(n20126), .B(n3032), .C(n24093), .CO(n20124), .S(n24091)
         );
  OR4X2 U23843 ( .A(n24068), .B(n24340), .C(n24308), .D(n24091), .Y(n20127) );
  OR4X2 U23844 ( .A(n24432), .B(n24389), .C(n24294), .D(n20127), .Y(n20128) );
  CMPR22X1 U23845 ( .A(n24300), .B(n20130), .CO(n20131), .S(n24301) );
  NOR2X1 U23846 ( .A(n20134), .B(n20133), .Y(n24066) );
  NOR2XL U23847 ( .A(n20137), .B(n24067), .Y(n20173) );
  OAI21XL U23848 ( .A0(n3030), .A1(n20140), .B0(n20139), .Y(n20211) );
  NAND3BX1 U23849 ( .AN(n20151), .B(n24722), .C(n20150), .Y(n20155) );
  NAND4BXL U23850 ( .AN(n20165), .B(n20164), .C(n24937), .D(n24938), .Y(n20166) );
  NAND2XL U23851 ( .A(n3030), .B(n20203), .Y(n20174) );
  OAI21XL U23852 ( .A0(n3030), .A1(n20175), .B0(n20174), .Y(n20212) );
  NAND2XL U23853 ( .A(n20213), .B(n3032), .Y(n20180) );
  OAI21XL U23854 ( .A0(n20212), .A1(n20138), .B0(n20180), .Y(n20244) );
  OAI22XL U23855 ( .A0(n3069), .A1(n20181), .B0(n20244), .B1(n20182), .Y(
        n20210) );
  NOR2XL U23856 ( .A(n20210), .B(n3075), .Y(n20193) );
  NAND2XL U23857 ( .A(n3030), .B(n20254), .Y(n20183) );
  OAI21XL U23858 ( .A0(n3030), .A1(n20092), .B0(n20183), .Y(n24719) );
  NAND2XL U23859 ( .A(n3030), .B(n20235), .Y(n20184) );
  OAI21XL U23860 ( .A0(n3030), .A1(n20185), .B0(n20184), .Y(n20250) );
  OAI22XL U23861 ( .A0(n3072), .A1(n24719), .B0(n20250), .B1(n3032), .Y(n24801) );
  NAND2XL U23862 ( .A(n3030), .B(n20195), .Y(n20187) );
  OAI21XL U23863 ( .A0(n3030), .A1(n20219), .B0(n20187), .Y(n20215) );
  NOR2XL U23864 ( .A(n3030), .B(n20088), .Y(n20190) );
  NAND2XL U23865 ( .A(n20248), .B(n3032), .Y(n20191) );
  OAI21XL U23866 ( .A0(n20215), .A1(n3032), .B0(n20191), .Y(n20245) );
  OAI22XL U23867 ( .A0(n20182), .A1(n24801), .B0(n20245), .B1(n3069), .Y(
        n24947) );
  NOR2XL U23868 ( .A(n24947), .B(n20066), .Y(n20192) );
  NAND2XL U23869 ( .A(n3030), .B(n20196), .Y(n20197) );
  OAI21XL U23870 ( .A0(n3030), .A1(n20198), .B0(n20197), .Y(n20217) );
  NAND2XL U23871 ( .A(n3030), .B(n20199), .Y(n20200) );
  OAI21XL U23872 ( .A0(n3030), .A1(n20201), .B0(n20200), .Y(n20224) );
  OAI22XL U23873 ( .A0(n3072), .A1(n20217), .B0(n20224), .B1(n3032), .Y(n20241) );
  NOR2XL U23874 ( .A(n20202), .B(n20138), .Y(n20208) );
  NAND2XL U23875 ( .A(n3030), .B(n20204), .Y(n20205) );
  OAI21XL U23876 ( .A0(n3030), .A1(n20206), .B0(n20205), .Y(n20223) );
  NOR2XL U23877 ( .A(n20223), .B(n3072), .Y(n20207) );
  OAI21XL U23878 ( .A0(n24894), .A1(n20241), .B0(n20209), .Y(n24684) );
  NAND2XL U23879 ( .A(n20210), .B(n3075), .Y(n24949) );
  NOR2XL U23880 ( .A(n24949), .B(n23200), .Y(n20996) );
  OAI22XL U23881 ( .A0(n3072), .A1(n20212), .B0(n20211), .B1(n20138), .Y(
        n20229) );
  NAND2XL U23882 ( .A(n20213), .B(n3072), .Y(n20214) );
  OAI21XL U23883 ( .A0(n3072), .A1(n20215), .B0(n20214), .Y(n20251) );
  OAI22XL U23884 ( .A0(n24721), .A1(n20066), .B0(n20216), .B1(n3075), .Y(
        n25352) );
  INVXL U23885 ( .A(n20217), .Y(n20222) );
  NOR2XL U23886 ( .A(n3030), .B(n20218), .Y(n20221) );
  AOI22XL U23887 ( .A0(n20222), .A1(n3072), .B0(n20239), .B1(n3032), .Y(n20259) );
  OAI22XL U23888 ( .A0(n3072), .A1(n20224), .B0(n20223), .B1(n3032), .Y(n20231) );
  OAI21XL U23889 ( .A0(n20225), .A1(n3075), .B0(n3074), .Y(n20226) );
  NAND2XL U23890 ( .A(n24570), .B(n24577), .Y(n20227) );
  OAI22XL U23891 ( .A0(n20229), .A1(n24894), .B0(n3069), .B1(n20228), .Y(
        n20252) );
  OAI22XL U23892 ( .A0(n20231), .A1(n24894), .B0(n20230), .B1(n3069), .Y(
        n20260) );
  NAND2XL U23893 ( .A(n20260), .B(n3075), .Y(n24902) );
  NOR2XL U23894 ( .A(n24902), .B(n23200), .Y(n24497) );
  NAND2XL U23895 ( .A(n24492), .B(n24497), .Y(n20233) );
  NOR2XL U23896 ( .A(n24835), .B(n23200), .Y(n20683) );
  NAND2XL U23897 ( .A(n20683), .B(n24462), .Y(n24476) );
  NAND2XL U23898 ( .A(n3030), .B(n20236), .Y(n20237) );
  OAI21XL U23899 ( .A0(n3030), .A1(n20238), .B0(n20237), .Y(n20258) );
  NAND2XL U23900 ( .A(n20239), .B(n3072), .Y(n20240) );
  OAI22XL U23901 ( .A0(n20241), .A1(n3069), .B0(n24683), .B1(n24894), .Y(
        n24833) );
  OAI22XL U23902 ( .A0(n20182), .A1(n20245), .B0(n20244), .B1(n3069), .Y(
        n24797) );
  NAND2XL U23903 ( .A(n24611), .B(n24607), .Y(n24646) );
  NAND2XL U23904 ( .A(n20248), .B(n3072), .Y(n20249) );
  OAI21XL U23905 ( .A0(n3072), .A1(n20250), .B0(n20249), .Y(n24720) );
  OAI22XL U23906 ( .A0(n20182), .A1(n24720), .B0(n20251), .B1(n3069), .Y(
        n24848) );
  NAND2XL U23907 ( .A(n3030), .B(n20255), .Y(n20256) );
  OAI21XL U23908 ( .A0(n3030), .A1(n20257), .B0(n20256), .Y(n24681) );
  OAI22XL U23909 ( .A0(n3072), .A1(n24681), .B0(n20258), .B1(n3032), .Y(n24751) );
  NOR2XL U23910 ( .A(n20260), .B(n3075), .Y(n20261) );
  AOI21XL U23911 ( .A0(n24898), .A1(n3075), .B0(n20261), .Y(n24651) );
  NAND2XL U23912 ( .A(n24630), .B(n24651), .Y(n20262) );
  NAND2XL U23913 ( .A(n24760), .B(n24811), .Y(n20263) );
  AOI22XL U23914 ( .A0(n25485), .A1(n3025), .B0(n24958), .B1(y11[12]), .Y(
        n20266) );
  NAND2XL U23915 ( .A(n20610), .B(n20706), .Y(n20271) );
  NOR2X1 U23916 ( .A(n20810), .B(n20271), .Y(n20272) );
  XOR2X2 U23917 ( .A(n20274), .B(n20704), .Y(n20615) );
  AOI22XL U23918 ( .A0(n20627), .A1(n23949), .B0(n23940), .B1(n23947), .Y(
        n20300) );
  INVXL U23919 ( .A(n20666), .Y(n20302) );
  NOR2XL U23920 ( .A(n23709), .B(n20302), .Y(n20303) );
  NOR2XL U23921 ( .A(n23709), .B(n23648), .Y(n20304) );
  XOR2X1 U23922 ( .A(n20306), .B(n20305), .Y(n23793) );
  AOI22X1 U23923 ( .A0(n3081), .A1(n23702), .B0(n23793), .B1(n4267), .Y(n24744) );
  INVXL U23924 ( .A(n20670), .Y(n20307) );
  NAND2XL U23925 ( .A(n3895), .B(n20308), .Y(n20310) );
  XOR2X1 U23926 ( .A(n20310), .B(n20309), .Y(n24220) );
  NOR2X4 U23927 ( .A(n5985), .B(n3121), .Y(n23794) );
  NAND2XL U23928 ( .A(n24211), .B(n23795), .Y(n20313) );
  INVXL U23929 ( .A(n20317), .Y(n20318) );
  XNOR2X1 U23930 ( .A(n3895), .B(n20318), .Y(n25298) );
  OAI21XL U23931 ( .A0(n3045), .A1(n25900), .B0(n20319), .Y(n20320) );
  INVXL U23932 ( .A(n20967), .Y(n20322) );
  NOR2XL U23933 ( .A(n20322), .B(n20326), .Y(n20323) );
  INVXL U23934 ( .A(n20333), .Y(n20334) );
  NAND2XL U23935 ( .A(n3357), .B(n20334), .Y(n20336) );
  NAND2X1 U23936 ( .A(n20337), .B(n5336), .Y(n20338) );
  NOR2X2 U23937 ( .A(n25813), .B(n3120), .Y(n25785) );
  XOR2X1 U23938 ( .A(n20342), .B(n20341), .Y(n20747) );
  NAND2X1 U23939 ( .A(n20343), .B(n5336), .Y(n20344) );
  NAND2XL U23940 ( .A(n3956), .B(n20348), .Y(n20349) );
  NOR2XL U23941 ( .A(n20929), .B(n20349), .Y(n20350) );
  NAND2XL U23942 ( .A(n3357), .B(n20356), .Y(n20357) );
  NAND2XL U23943 ( .A(n20363), .B(n20618), .Y(n20364) );
  OR2XL U23944 ( .A(n3024), .B(valid[0]), .Y(n20860) );
  NOR2XL U23945 ( .A(n20376), .B(n20375), .Y(n23189) );
  NOR2XL U23946 ( .A(n20377), .B(n23189), .Y(n20383) );
  OAI21XL U23947 ( .A0(n3067), .A1(n20387), .B0(n20386), .Y(n20481) );
  OAI21XL U23948 ( .A0(n3067), .A1(n20389), .B0(n20388), .Y(n20487) );
  OAI22XL U23949 ( .A0(n3031), .A1(n20481), .B0(n20487), .B1(n3071), .Y(n20504) );
  NOR2XL U23950 ( .A(n3067), .B(n20390), .Y(n20391) );
  AOI21XL U23951 ( .A0(n20443), .A1(n3067), .B0(n20391), .Y(n20489) );
  NOR2XL U23952 ( .A(n20392), .B(n3071), .Y(n20393) );
  NAND2XL U23953 ( .A(n20506), .B(n20473), .Y(n20394) );
  OAI21XL U23954 ( .A0(n20473), .A1(n20504), .B0(n20394), .Y(n20427) );
  OAI22XL U23955 ( .A0(n20427), .A1(n20597), .B0(n20395), .B1(n20576), .Y(
        n20519) );
  OAI21XL U23956 ( .A0(n3067), .A1(n20397), .B0(n20396), .Y(n20594) );
  OAI21XL U23957 ( .A0(n3067), .A1(n20399), .B0(n20398), .Y(n20531) );
  OAI22XL U23958 ( .A0(n3031), .A1(n20594), .B0(n20531), .B1(n3071), .Y(n20553) );
  AOI21XL U23959 ( .A0(n20561), .A1(n3067), .B0(n20401), .Y(n20592) );
  OAI21XL U23960 ( .A0(n3067), .A1(n20403), .B0(n3071), .Y(n20406) );
  AOI21XL U23961 ( .A0(n3031), .A1(n20592), .B0(n20407), .Y(n20408) );
  OAI21XL U23962 ( .A0(n3068), .A1(n20553), .B0(n20409), .Y(n20423) );
  NOR2XL U23963 ( .A(n3067), .B(n20410), .Y(n20413) );
  NOR2XL U23964 ( .A(n3067), .B(n20414), .Y(n20417) );
  AOI22XL U23965 ( .A0(n20482), .A1(n3031), .B0(n20484), .B1(n3071), .Y(n20505) );
  OAI21XL U23966 ( .A0(n3067), .A1(n20419), .B0(n20418), .Y(n20530) );
  OAI21XL U23967 ( .A0(n3067), .A1(n20421), .B0(n20420), .Y(n20486) );
  OAI22XL U23968 ( .A0(n3031), .A1(n20530), .B0(n20486), .B1(n3071), .Y(n20555) );
  NAND2XL U23969 ( .A(n20426), .B(n20576), .Y(n20429) );
  NAND2XL U23970 ( .A(n3067), .B(n20432), .Y(n20433) );
  OAI21XL U23971 ( .A0(n3067), .A1(n20434), .B0(n20433), .Y(n20471) );
  OAI21XL U23972 ( .A0(n3067), .A1(n20438), .B0(n20437), .Y(n20475) );
  OAI22XL U23973 ( .A0(n3031), .A1(n20471), .B0(n20475), .B1(n3071), .Y(n20510) );
  INVXL U23974 ( .A(n20439), .Y(n20442) );
  NAND2XL U23975 ( .A(n3067), .B(n20440), .Y(n20441) );
  OAI21XL U23976 ( .A0(n3067), .A1(n20442), .B0(n20441), .Y(n20474) );
  NOR2XL U23977 ( .A(n3067), .B(n20444), .Y(n20447) );
  NAND2XL U23978 ( .A(n20476), .B(n3031), .Y(n20448) );
  OAI21XL U23979 ( .A0(n3031), .A1(n20474), .B0(n20448), .Y(n20513) );
  OAI22XL U23980 ( .A0(n20473), .A1(n20510), .B0(n20513), .B1(n3068), .Y(
        n20522) );
  NOR2XL U23981 ( .A(n20522), .B(n20576), .Y(n20468) );
  NAND2XL U23982 ( .A(n3067), .B(n20450), .Y(n20451) );
  OAI21XL U23983 ( .A0(n3067), .A1(n20452), .B0(n20451), .Y(n20546) );
  OAI21XL U23984 ( .A0(n3067), .A1(n20456), .B0(n20455), .Y(n20470) );
  OAI22XL U23985 ( .A0(n3031), .A1(n20546), .B0(n20470), .B1(n3071), .Y(n20568) );
  NAND2XL U23986 ( .A(n3067), .B(n20458), .Y(n20459) );
  OAI21XL U23987 ( .A0(n3067), .A1(n20460), .B0(n20459), .Y(n20469) );
  NAND2XL U23988 ( .A(n3067), .B(n20461), .Y(n20462) );
  OAI21XL U23989 ( .A0(n3067), .A1(n20463), .B0(n20462), .Y(n20472) );
  OAI22XL U23990 ( .A0(n3031), .A1(n20469), .B0(n20472), .B1(n3071), .Y(n20511) );
  NOR2XL U23991 ( .A(n20511), .B(n3068), .Y(n20464) );
  OAI22XL U23992 ( .A0(n20468), .A1(n20467), .B0(n20466), .B1(n3073), .Y(
        n24793) );
  NAND2XL U23993 ( .A(n24785), .B(n4779), .Y(n20493) );
  OAI22XL U23994 ( .A0(n3031), .A1(n20470), .B0(n20469), .B1(n3071), .Y(n20541) );
  OAI22XL U23995 ( .A0(n3031), .A1(n20472), .B0(n20471), .B1(n3071), .Y(n20495) );
  OAI22XL U23996 ( .A0(n20473), .A1(n20541), .B0(n20495), .B1(n3068), .Y(
        n20577) );
  OAI22XL U23997 ( .A0(n3031), .A1(n20475), .B0(n20474), .B1(n3071), .Y(n20494) );
  AOI22XL U23998 ( .A0(n20477), .A1(n3031), .B0(n20476), .B1(n3071), .Y(n20496) );
  NAND2XL U23999 ( .A(n20496), .B(n20473), .Y(n20478) );
  NOR2XL U24000 ( .A(n20517), .B(n20576), .Y(n20479) );
  INVXL U24001 ( .A(n20481), .Y(n20483) );
  AOI22XL U24002 ( .A0(n20483), .A1(n3031), .B0(n20482), .B1(n3071), .Y(n20499) );
  NAND2XL U24003 ( .A(n20484), .B(n3031), .Y(n20485) );
  OAI21XL U24004 ( .A0(n3031), .A1(n20486), .B0(n20485), .Y(n20535) );
  NOR2XL U24005 ( .A(n20487), .B(n3031), .Y(n20488) );
  AOI21XL U24006 ( .A0(n20489), .A1(n3031), .B0(n20488), .Y(n20501) );
  NAND2XL U24007 ( .A(n20501), .B(n3068), .Y(n20490) );
  OAI21XL U24008 ( .A0(n3068), .A1(n20491), .B0(n20490), .Y(n20518) );
  NOR2XL U24009 ( .A(n20518), .B(n20576), .Y(n20492) );
  AOI21XL U24010 ( .A0(n20598), .A1(n20576), .B0(n20492), .Y(n20841) );
  NAND2XL U24011 ( .A(n24712), .B(n20841), .Y(n24784) );
  OAI22XL U24012 ( .A0(n20473), .A1(n20495), .B0(n20494), .B1(n3068), .Y(
        n20550) );
  NOR2XL U24013 ( .A(n20526), .B(n20576), .Y(n20497) );
  NAND2XL U24014 ( .A(n20499), .B(n3068), .Y(n20500) );
  NAND2XL U24015 ( .A(n20506), .B(n3068), .Y(n20507) );
  NOR2XL U24016 ( .A(n20524), .B(n20576), .Y(n20509) );
  OAI22XL U24017 ( .A0(n20473), .A1(n20511), .B0(n20510), .B1(n3068), .Y(
        n20572) );
  OAI22XL U24018 ( .A0(n20513), .A1(n20473), .B0(n20512), .B1(n3068), .Y(
        n20525) );
  NAND2XL U24019 ( .A(n20906), .B(n20877), .Y(n20515) );
  NAND2XL U24020 ( .A(n20518), .B(n20576), .Y(n20602) );
  OAI21XL U24021 ( .A0(n20520), .A1(n20576), .B0(n3073), .Y(n20521) );
  NAND2XL U24022 ( .A(n24566), .B(n20889), .Y(n20523) );
  NAND2XL U24023 ( .A(n20524), .B(n20576), .Y(n20560) );
  NAND2XL U24024 ( .A(n20525), .B(n20576), .Y(n20574) );
  NAND2XL U24025 ( .A(n20918), .B(n20913), .Y(n20527) );
  NAND2XL U24026 ( .A(n20526), .B(n20576), .Y(n20552) );
  NAND2XL U24027 ( .A(n23773), .B(n25301), .Y(n20909) );
  NOR2X2 U24028 ( .A(n20529), .B(n20838), .Y(n23829) );
  NOR2XL U24029 ( .A(n20530), .B(n3071), .Y(n20533) );
  NOR2XL U24030 ( .A(n20531), .B(n3031), .Y(n20532) );
  AOI21XL U24031 ( .A0(n20591), .A1(n3068), .B0(n20597), .Y(n20534) );
  OAI21XL U24032 ( .A0(n3068), .A1(n20535), .B0(n20534), .Y(n20536) );
  INVXL U24033 ( .A(n20536), .Y(n20540) );
  NOR2XL U24034 ( .A(n20537), .B(n20576), .Y(n20539) );
  NOR2XL U24035 ( .A(n20541), .B(n3068), .Y(n20548) );
  NAND2XL U24036 ( .A(n3067), .B(n20543), .Y(n20544) );
  OAI21XL U24037 ( .A0(n3067), .A1(n20545), .B0(n20544), .Y(n20565) );
  OAI22XL U24038 ( .A0(n3031), .A1(n20565), .B0(n20546), .B1(n3071), .Y(n20578) );
  OAI21XL U24039 ( .A0(n20578), .A1(n20473), .B0(n20576), .Y(n20547) );
  OAI21XL U24040 ( .A0(n20576), .A1(n20550), .B0(n20549), .Y(n20551) );
  OAI21XL U24041 ( .A0(n20552), .A1(n3073), .B0(n20551), .Y(n23608) );
  NAND2XL U24042 ( .A(n23754), .B(n23608), .Y(n23827) );
  OAI21XL U24043 ( .A0(n3068), .A1(n20555), .B0(n20554), .Y(n20558) );
  NAND2XL U24044 ( .A(n20556), .B(n20597), .Y(n20557) );
  OAI21XL U24045 ( .A0(n20560), .A1(n3073), .B0(n20559), .Y(n23616) );
  OAI21XL U24046 ( .A0(n3067), .A1(n20564), .B0(n20563), .Y(n20583) );
  OAI21XL U24047 ( .A0(n20583), .A1(n3031), .B0(n3068), .Y(n20567) );
  NOR2XL U24048 ( .A(n20565), .B(n3071), .Y(n20566) );
  OAI21XL U24049 ( .A0(n20567), .A1(n20566), .B0(n20576), .Y(n20570) );
  NOR2XL U24050 ( .A(n20568), .B(n3068), .Y(n20569) );
  OAI21XL U24051 ( .A0(n20572), .A1(n20576), .B0(n20571), .Y(n20573) );
  NAND2XL U24052 ( .A(n23616), .B(n23833), .Y(n20575) );
  NOR2XL U24053 ( .A(n20577), .B(n20576), .Y(n20589) );
  NOR2XL U24054 ( .A(n20578), .B(n3068), .Y(n20587) );
  OAI21XL U24055 ( .A0(n20585), .A1(n20584), .B0(n20576), .Y(n20586) );
  NAND2XL U24056 ( .A(n20591), .B(n20473), .Y(n20596) );
  OAI21XL U24057 ( .A0(n3071), .A1(n20594), .B0(n20593), .Y(n20595) );
  NAND2XL U24058 ( .A(n20598), .B(n20597), .Y(n20599) );
  NAND2XL U24059 ( .A(n23829), .B(n20604), .Y(n20606) );
  XOR2X1 U24060 ( .A(n20606), .B(n20605), .Y(n20607) );
  AOI222X1 U24061 ( .A0(n25828), .A1(n25737), .B0(n25743), .B1(y20[22]), .C0(
        n25824), .C1(n20890), .Y(n2382) );
  NOR2XL U24062 ( .A(n20609), .B(n20704), .Y(n20611) );
  NAND2XL U24063 ( .A(n20611), .B(n20610), .Y(n20612) );
  NAND2XL U24064 ( .A(n23829), .B(n23798), .Y(n20633) );
  XOR2X1 U24065 ( .A(n20633), .B(n23799), .Y(n20634) );
  INVXL U24066 ( .A(n20790), .Y(n20645) );
  NOR2X1 U24067 ( .A(n20647), .B(n20646), .Y(n20648) );
  AOI22XL U24068 ( .A0(n20659), .A1(n25807), .B0(n2983), .B1(temp2[23]), .Y(
        n20660) );
  NAND2XL U24069 ( .A(n23744), .B(n20662), .Y(n20664) );
  NAND2XL U24070 ( .A(n20666), .B(n20665), .Y(n20667) );
  XOR2X1 U24071 ( .A(n20673), .B(n20672), .Y(n24227) );
  NAND2XL U24072 ( .A(n24227), .B(n23795), .Y(n20674) );
  INVXL U24073 ( .A(n20677), .Y(n20679) );
  NAND2XL U24074 ( .A(n20679), .B(n20678), .Y(n20680) );
  XOR2X1 U24075 ( .A(n23482), .B(n20680), .Y(n23483) );
  INVXL U24076 ( .A(n20683), .Y(n20681) );
  XNOR2XL U24077 ( .A(n20681), .B(n24462), .Y(n20682) );
  AOI22XL U24078 ( .A0(n25623), .A1(n3025), .B0(n24958), .B1(y11[1]), .Y(
        n20685) );
  INVXL U24079 ( .A(n3009), .Y(n20694) );
  NAND2XL U24080 ( .A(n20694), .B(n20693), .Y(n20695) );
  AOI22X1 U24081 ( .A0(n21051), .A1(n5336), .B0(n3136), .B1(n24263), .Y(n25293) );
  INVXL U24082 ( .A(n4651), .Y(n20702) );
  NOR2X1 U24083 ( .A(n20708), .B(n20707), .Y(n20710) );
  AOI22XL U24084 ( .A0(n25727), .A1(n25724), .B0(n25723), .B1(temp0[22]), .Y(
        n20729) );
  INVXL U24085 ( .A(n20735), .Y(n20737) );
  NOR2XL U24086 ( .A(n20737), .B(n20736), .Y(n20738) );
  INVXL U24087 ( .A(n20750), .Y(n2302) );
  NAND2X1 U24088 ( .A(n3132), .B(n20751), .Y(n20753) );
  NOR2XL U24089 ( .A(n20760), .B(n20845), .Y(n20761) );
  XOR2X1 U24090 ( .A(n20764), .B(n20763), .Y(n20847) );
  AOI22XL U24091 ( .A0(n20824), .A1(n23949), .B0(n23933), .B1(n23947), .Y(
        n20773) );
  AND2X2 U24092 ( .A(n25128), .B(n20795), .Y(n20777) );
  INVXL U24093 ( .A(n25176), .Y(n20785) );
  INVXL U24094 ( .A(n20780), .Y(n20781) );
  INVXL U24095 ( .A(n20791), .Y(n20789) );
  AOI2BB2X1 U24096 ( .B0(n2984), .B1(temp2[24]), .A0N(n25709), .A1N(n4582), 
        .Y(n20793) );
  AND2X2 U24097 ( .A(n25128), .B(n25124), .Y(n20796) );
  AOI211X1 U24098 ( .A0(n5911), .A1(n20797), .B0(n20796), .C0(n25127), .Y(
        n25207) );
  INVXL U24099 ( .A(n25207), .Y(n20806) );
  ADDHXL U24100 ( .A(n20800), .B(n20799), .CO(n24268), .S(n20780) );
  AOI2BB2XL U24101 ( .B0(n2984), .B1(temp2[29]), .A0N(n25842), .A1N(n4581), 
        .Y(n20805) );
  OAI2BB1XL U24102 ( .A0N(n25807), .A1N(n20806), .B0(n20805), .Y(n2559) );
  NAND2XL U24103 ( .A(n20808), .B(n20807), .Y(n20809) );
  NOR2XL U24104 ( .A(n20810), .B(n20809), .Y(n20811) );
  AOI22XL U24105 ( .A0(n23544), .A1(n23949), .B0(n23947), .B1(n20824), .Y(
        n20825) );
  INVXL U24106 ( .A(n20828), .Y(n20829) );
  NAND2XL U24107 ( .A(n20829), .B(n20865), .Y(n20834) );
  INVXL U24108 ( .A(n20830), .Y(n20836) );
  NOR2XL U24109 ( .A(n20834), .B(n20836), .Y(n20831) );
  XOR2X1 U24110 ( .A(n20833), .B(n3148), .Y(n23893) );
  INVXL U24111 ( .A(n20834), .Y(n20835) );
  NAND2X1 U24112 ( .A(n5100), .B(n20835), .Y(n20837) );
  XOR2X1 U24113 ( .A(n20837), .B(n20836), .Y(n20872) );
  NAND2XL U24114 ( .A(n24789), .B(n20848), .Y(n20839) );
  XOR2X1 U24115 ( .A(n20839), .B(n24707), .Y(n20840) );
  AOI222X1 U24116 ( .A0(n24677), .A1(n25737), .B0(n25743), .B1(y20[12]), .C0(
        n25486), .C1(n20890), .Y(n2372) );
  OAI21XL U24117 ( .A0(n3045), .A1(n25913), .B0(n20842), .Y(n20843) );
  NAND2X1 U24118 ( .A(n5100), .B(n3586), .Y(n20846) );
  XOR2X1 U24119 ( .A(n20846), .B(n20845), .Y(n23894) );
  INVXL U24120 ( .A(n20848), .Y(n24787) );
  NOR2XL U24121 ( .A(n24787), .B(n24784), .Y(n20849) );
  NAND2XL U24122 ( .A(n20849), .B(n24789), .Y(n20851) );
  INVXL U24123 ( .A(n24785), .Y(n20850) );
  AOI222X1 U24124 ( .A0(n24743), .A1(n25737), .B0(n25743), .B1(y20[14]), .C0(
        n25460), .C1(n20890), .Y(n2374) );
  NAND2XL U24125 ( .A(n5100), .B(n20865), .Y(n20854) );
  NAND2XL U24126 ( .A(n20856), .B(n20855), .Y(n20878) );
  NOR2XL U24127 ( .A(n20878), .B(n20880), .Y(n20857) );
  CLKINVX3 U24128 ( .A(n20860), .Y(n25744) );
  NAND2XL U24129 ( .A(n24789), .B(n23583), .Y(n20862) );
  INVXL U24130 ( .A(n20864), .Y(n20861) );
  XOR2X1 U24131 ( .A(n20862), .B(n20861), .Y(n20863) );
  AOI222X1 U24132 ( .A0(n23579), .A1(n25744), .B0(n25743), .B1(y20[9]), .C0(
        n25520), .C1(n20890), .Y(n2369) );
  INVXL U24133 ( .A(n20865), .Y(n20867) );
  NOR2XL U24134 ( .A(n20867), .B(n20866), .Y(n20868) );
  NOR2XL U24135 ( .A(n20901), .B(n20903), .Y(n20873) );
  NAND2XL U24136 ( .A(n24789), .B(n20873), .Y(n20875) );
  AOI222X1 U24137 ( .A0(n23658), .A1(n25744), .B0(n25743), .B1(y20[11]), .C0(
        n25496), .C1(n20890), .Y(n2371) );
  INVXL U24138 ( .A(n20878), .Y(n20879) );
  NAND2XL U24139 ( .A(n5125), .B(n20879), .Y(n20881) );
  INVXL U24140 ( .A(n24561), .Y(n20883) );
  NAND2XL U24141 ( .A(n20883), .B(n24566), .Y(n20885) );
  NOR2XL U24142 ( .A(n20885), .B(n24562), .Y(n20887) );
  INVXL U24143 ( .A(n20889), .Y(n20886) );
  INVXL U24144 ( .A(n20894), .Y(n20891) );
  INVXL U24145 ( .A(n20898), .Y(n23621) );
  AOI222X1 U24146 ( .A0(n24526), .A1(n25744), .B0(n25743), .B1(y20[4]), .C0(
        n25578), .C1(n20890), .Y(n2364) );
  INVXL U24147 ( .A(n20901), .Y(n20902) );
  NAND2XL U24148 ( .A(n24789), .B(n20902), .Y(n20904) );
  INVXL U24149 ( .A(n20909), .Y(n20916) );
  NAND2XL U24150 ( .A(n20916), .B(n20918), .Y(n20911) );
  INVXL U24151 ( .A(n20913), .Y(n20910) );
  AOI22X1 U24152 ( .A0(n20385), .A1(n20913), .B0(n25300), .B1(n20912), .Y(
        n24512) );
  INVXL U24153 ( .A(n20918), .Y(n20915) );
  AOI222X1 U24154 ( .A0(n24490), .A1(n25744), .B0(n25743), .B1(y20[2]), .C0(
        n25610), .C1(n20890), .Y(n2362) );
  NAND2XL U24155 ( .A(n20927), .B(n20920), .Y(n20921) );
  INVXL U24156 ( .A(n20941), .Y(n2338) );
  AOI22XL U24157 ( .A0(n23949), .A1(n20962), .B0(n23947), .B1(n20961), .Y(
        n20963) );
  INVXL U24158 ( .A(n20966), .Y(n20968) );
  NAND2XL U24159 ( .A(n20968), .B(n20967), .Y(n21031) );
  INVXL U24160 ( .A(n21031), .Y(n20969) );
  INVX1 U24161 ( .A(n20970), .Y(n21030) );
  INVXL U24162 ( .A(n20972), .Y(n20973) );
  OR2X2 U24163 ( .A(n24145), .B(n4581), .Y(n20977) );
  NAND3X1 U24164 ( .A(n20979), .B(n20978), .C(n20977), .Y(n2547) );
  INVXL U24165 ( .A(n20980), .Y(n20985) );
  NOR2XL U24166 ( .A(n20985), .B(n20983), .Y(n20981) );
  INVXL U24167 ( .A(n20990), .Y(n20991) );
  AOI22XL U24168 ( .A0(n25577), .A1(n3025), .B0(n24958), .B1(y11[4]), .Y(
        n20998) );
  OAI21XL U24169 ( .A0(n25271), .A1(n21002), .B0(n21001), .Y(n24918) );
  NAND2XL U24170 ( .A(n21003), .B(n3127), .Y(n21004) );
  OAI21XL U24171 ( .A0(n3127), .A1(n24918), .B0(n21004), .Y(n25015) );
  OAI21XL U24172 ( .A0(n25015), .A1(n15808), .B0(n3077), .Y(n21007) );
  NOR2XL U24173 ( .A(n21005), .B(n3125), .Y(n21006) );
  NOR2XL U24174 ( .A(n21008), .B(n3077), .Y(n21010) );
  NAND2XL U24175 ( .A(n25286), .B(n4782), .Y(n21013) );
  OAI21XL U24176 ( .A0(n25059), .A1(n25921), .B0(n21015), .Y(n21016) );
  NOR2XL U24177 ( .A(n21022), .B(n21024), .Y(n21018) );
  INVXL U24178 ( .A(n21022), .Y(n21023) );
  OAI21XL U24179 ( .A0(n3045), .A1(n25903), .B0(n21025), .Y(n21026) );
  OAI21XL U24180 ( .A0(n3045), .A1(n25906), .B0(n21027), .Y(n21028) );
  NOR2XL U24181 ( .A(n21031), .B(n21030), .Y(n21032) );
  OAI21XL U24182 ( .A0(n3045), .A1(n25904), .B0(n21033), .Y(n21034) );
  NOR2XL U24183 ( .A(n5410), .B(n21037), .Y(n21038) );
  NAND2XL U24184 ( .A(n3895), .B(n21038), .Y(n21040) );
  XOR2X1 U24185 ( .A(n21040), .B(n21039), .Y(n24174) );
  OAI21XL U24186 ( .A0(n3045), .A1(n26234), .B0(n21041), .Y(n21042) );
  NAND2XL U24187 ( .A(n5978), .B(n21043), .Y(n21044) );
  OAI21XL U24188 ( .A0(n3045), .A1(n25914), .B0(n21046), .Y(n21047) );
  AOI22X1 U24189 ( .A0(n21052), .A1(n5336), .B0(n3136), .B1(n21051), .Y(n24116) );
  NOR2X4 U24190 ( .A(n21057), .B(n21056), .Y(n23152) );
  OAI21XL U24191 ( .A0(n11089), .A1(n22989), .B0(n4707), .Y(M6_mult_x_15_n634)
         );
  INVX1 U24192 ( .A(n22990), .Y(n22737) );
  AND3X2 U24193 ( .A(n21072), .B(n21071), .C(n21070), .Y(n22927) );
  OAI21XL U24194 ( .A0(n22913), .A1(n22909), .B0(n21060), .Y(n21061) );
  AND3X2 U24195 ( .A(n22563), .B(n22562), .C(n21064), .Y(n22976) );
  OAI21XL U24196 ( .A0(n11082), .A1(n22984), .B0(n21065), .Y(n21066) );
  NOR2X4 U24197 ( .A(n21072), .B(n21071), .Y(n22928) );
  OAI21XL U24198 ( .A0(n23076), .A1(n22909), .B0(n21074), .Y(n21075) );
  OAI21XL U24199 ( .A0(n22924), .A1(n22909), .B0(n21076), .Y(n21077) );
  INVX1 U24200 ( .A(n22713), .Y(n26489) );
  NOR2X4 U24201 ( .A(n21082), .B(n21081), .Y(n23003) );
  AND3X2 U24202 ( .A(n21082), .B(n21081), .C(n21080), .Y(n23001) );
  AOI222XL U24203 ( .A0(n23003), .A1(n26496), .B0(n22969), .B1(n10775), .C0(
        n23001), .C1(n10769), .Y(n21083) );
  OAI21XL U24204 ( .A0(n22924), .A1(n23005), .B0(n21083), .Y(n21084) );
  XOR2XL U24205 ( .A(n21084), .B(n21089), .Y(M6_mult_x_15_n1129) );
  OAI21XL U24206 ( .A0(n23155), .A1(n23005), .B0(n21088), .Y(n21090) );
  NOR3XL U24207 ( .A(iter[2]), .B(iter[0]), .C(n26308), .Y(n21092) );
  NOR4BXL U24208 ( .AN(n26309), .B(iter[1]), .C(iter[5]), .D(iter[6]), .Y(
        n21091) );
  NAND4XL U24209 ( .A(iter[4]), .B(iter[8]), .C(n21092), .D(n21091), .Y(n21100) );
  NAND2X1 U24210 ( .A(n23997), .B(n21100), .Y(n25856) );
  NAND2XL U24211 ( .A(n2972), .B(iter[0]), .Y(n23063) );
  INVXL U24212 ( .A(learning_rate[26]), .Y(n21104) );
  NOR2XL U24213 ( .A(learning_rate[23]), .B(learning_rate[24]), .Y(n24003) );
  NAND2XL U24214 ( .A(n24003), .B(n24006), .Y(n24002) );
  NOR2XL U24215 ( .A(n24002), .B(learning_rate[26]), .Y(n23051) );
  AOI21XL U24216 ( .A0(n24002), .A1(learning_rate[26]), .B0(n23051), .Y(n21102) );
  NAND4XL U24217 ( .A(learning_rate[23]), .B(learning_rate[24]), .C(
        learning_rate[25]), .D(learning_rate[26]), .Y(n21094) );
  NOR2XL U24218 ( .A(n21094), .B(n23053), .Y(n21099) );
  NAND2XL U24219 ( .A(n21099), .B(learning_rate[28]), .Y(n21098) );
  NOR2XL U24220 ( .A(n21098), .B(n21093), .Y(n21101) );
  OR2XL U24221 ( .A(n21101), .B(learning_rate[30]), .Y(n23976) );
  AOI21XL U24222 ( .A0(n21098), .A1(n21093), .B0(n21101), .Y(n23977) );
  INVXL U24223 ( .A(n21099), .Y(n21097) );
  NAND2XL U24224 ( .A(n21094), .B(n23053), .Y(n21096) );
  NOR2BXL U24225 ( .AN(n21094), .B(n23051), .Y(n21095) );
  AOI21XL U24226 ( .A0(n21097), .A1(n21096), .B0(n21095), .Y(n21106) );
  OAI21XL U24227 ( .A0(n21099), .A1(learning_rate[28]), .B0(n21098), .Y(n21105) );
  NAND2XL U24228 ( .A(n21106), .B(n21105), .Y(n23978) );
  NOR2XL U24229 ( .A(n23977), .B(n23978), .Y(n24012) );
  INVXL U24230 ( .A(n24008), .Y(n22471) );
  NAND2XL U24231 ( .A(learning_rate[30]), .B(n21101), .Y(n24011) );
  AOI21XL U24232 ( .A0(n21104), .A1(n23985), .B0(n21103), .Y(n2625) );
  INVXL U24233 ( .A(learning_rate[28]), .Y(n21109) );
  OAI21XL U24234 ( .A0(n21106), .A1(n21105), .B0(n23978), .Y(n21107) );
  AOI21XL U24235 ( .A0(n24008), .A1(n21107), .B0(n24007), .Y(n21108) );
  AOI21XL U24236 ( .A0(n21109), .A1(n23985), .B0(n21108), .Y(n2623) );
  CMPR32X1 U24237 ( .A(n22698), .B(n23109), .C(n11073), .CO(M6_mult_x_15_n447), 
        .S(M6_mult_x_15_n448) );
  CMPR32X1 U24238 ( .A(n22967), .B(n23151), .C(n11059), .CO(M6_mult_x_15_n487), 
        .S(M6_mult_x_15_n488) );
  CLKINVX3 U24239 ( .A(n25848), .Y(n25428) );
  AOI21XL U24240 ( .A0(n25541), .A1(w1[361]), .B0(n21115), .Y(n1918) );
  AOI21XL U24241 ( .A0(n3216), .A1(w1[362]), .B0(n21117), .Y(n1922) );
  AOI21XL U24242 ( .A0(n25541), .A1(w1[229]), .B0(n21119), .Y(n1774) );
  AOI21XL U24243 ( .A0(n25541), .A1(w1[359]), .B0(n21121), .Y(n1910) );
  AOI21XL U24244 ( .A0(n25541), .A1(w1[360]), .B0(n21123), .Y(n1914) );
  OAI21XL U24245 ( .A0(n3117), .A1(n26348), .B0(n21124), .Y(n21125) );
  AOI21XL U24246 ( .A0(n25541), .A1(w1[231]), .B0(n21125), .Y(n1782) );
  OAI21XL U24247 ( .A0(n3117), .A1(n26347), .B0(n21126), .Y(n21127) );
  AOI21XL U24248 ( .A0(n25541), .A1(w1[232]), .B0(n21127), .Y(n1786) );
  OAI21XL U24249 ( .A0(n3117), .A1(n26346), .B0(n21128), .Y(n21129) );
  AOI21XL U24250 ( .A0(n25541), .A1(w1[233]), .B0(n21129), .Y(n1790) );
  AOI21XL U24251 ( .A0(n25541), .A1(w1[357]), .B0(n21131), .Y(n1902) );
  OAI21XL U24252 ( .A0(n3117), .A1(n26344), .B0(n21132), .Y(n21133) );
  AOI21XL U24253 ( .A0(n25541), .A1(w1[235]), .B0(n21133), .Y(n1798) );
  AOI21XL U24254 ( .A0(n25541), .A1(w1[364]), .B0(n21135), .Y(n1930) );
  OAI21XL U24255 ( .A0(n3117), .A1(n26343), .B0(n21136), .Y(n21137) );
  AOI21XL U24256 ( .A0(n25541), .A1(w1[236]), .B0(n21137), .Y(n1802) );
  OAI21XL U24257 ( .A0(n3117), .A1(n26337), .B0(n21138), .Y(n21139) );
  AOI21XL U24258 ( .A0(n25541), .A1(w1[244]), .B0(n21139), .Y(n1834) );
  OAI21XL U24259 ( .A0(n3117), .A1(n26336), .B0(n21140), .Y(n21141) );
  AOI21XL U24260 ( .A0(n25541), .A1(w1[245]), .B0(n21141), .Y(n1838) );
  OAI21XL U24261 ( .A0(n3117), .A1(n26334), .B0(n21142), .Y(n21143) );
  AOI21XL U24262 ( .A0(n25541), .A1(w1[248]), .B0(n21143), .Y(n1850) );
  OAI21XL U24263 ( .A0(n3117), .A1(n26335), .B0(n21144), .Y(n21145) );
  AOI21XL U24264 ( .A0(n25541), .A1(w1[255]), .B0(n21145), .Y(n1878) );
  AOI21XL U24265 ( .A0(n25541), .A1(w1[230]), .B0(n21147), .Y(n1778) );
  INVX8 U24266 ( .A(n3117), .Y(n25410) );
  AOI21XL U24267 ( .A0(n25541), .A1(w1[383]), .B0(n21149), .Y(n2006) );
  OAI21XL U24268 ( .A0(n3117), .A1(n26345), .B0(n21150), .Y(n21151) );
  AOI21XL U24269 ( .A0(n25541), .A1(w1[234]), .B0(n21151), .Y(n1794) );
  AOI21XL U24270 ( .A0(n25541), .A1(w1[358]), .B0(n21153), .Y(n1906) );
  AOI21XL U24271 ( .A0(n25541), .A1(w1[376]), .B0(n21155), .Y(n1978) );
  AOI21XL U24272 ( .A0(n25541), .A1(w1[246]), .B0(n21157), .Y(n1842) );
  AOI21XL U24273 ( .A0(n25541), .A1(w1[363]), .B0(n21159), .Y(n1926) );
  AOI21XL U24274 ( .A0(n25541), .A1(w1[373]), .B0(n21161), .Y(n1966) );
  AOI21XL U24275 ( .A0(n21112), .A1(w1[372]), .B0(n21163), .Y(n1962) );
  AOI21XL U24276 ( .A0(n25541), .A1(w1[374]), .B0(n21165), .Y(n1970) );
  AOI21XL U24277 ( .A0(w1[156]), .A1(n3028), .B0(n21172), .Y(n1994) );
  OAI21XL U24278 ( .A0(n6196), .A1(n21256), .B0(n21174), .Y(n21626) );
  OAI21XL U24279 ( .A0(n26140), .A1(n25887), .B0(w1[3]), .Y(n21176) );
  OAI21XL U24280 ( .A0(n26140), .A1(n25887), .B0(temp0[3]), .Y(n21178) );
  OAI21XL U24281 ( .A0(n26140), .A1(n25887), .B0(w1[1]), .Y(n21181) );
  NAND3XL U24282 ( .A(cs[0]), .B(cs[1]), .C(y20[1]), .Y(n21180) );
  OAI21XL U24283 ( .A0(n26140), .A1(n25887), .B0(temp0[1]), .Y(n21183) );
  OAI21XL U24284 ( .A0(n25887), .A1(n26140), .B0(w1[2]), .Y(n21186) );
  NAND3XL U24285 ( .A(cs[0]), .B(cs[1]), .C(y20[2]), .Y(n21185) );
  OAI21XL U24286 ( .A0(n26140), .A1(n25887), .B0(temp0[2]), .Y(n21188) );
  CLKINVX3 U24287 ( .A(n4631), .Y(n21311) );
  OAI21XL U24288 ( .A0(n6203), .A1(n21311), .B0(n21190), .Y(n21619) );
  OAI21XL U24289 ( .A0(n26140), .A1(n25887), .B0(w1[0]), .Y(n21192) );
  NAND3XL U24290 ( .A(cs[0]), .B(cs[1]), .C(y20[0]), .Y(n21191) );
  NAND2XL U24291 ( .A(n21619), .B(n21193), .Y(n21198) );
  OAI21XL U24292 ( .A0(n21199), .A1(n21198), .B0(n21197), .Y(n21206) );
  OAI21XL U24293 ( .A0(n21204), .A1(n21203), .B0(n21202), .Y(n21205) );
  INVX1 U24294 ( .A(n21530), .Y(n21225) );
  OAI21XL U24295 ( .A0(n6181), .A1(n21331), .B0(n21209), .Y(n21469) );
  OAI21XL U24296 ( .A0(n26181), .A1(n21256), .B0(n21210), .Y(n21600) );
  OAI21XL U24297 ( .A0(n6180), .A1(n21311), .B0(n21211), .Y(n21556) );
  OAI21XL U24298 ( .A0(n6214), .A1(n21256), .B0(n21214), .Y(n21554) );
  OAI21XL U24299 ( .A0(n26183), .A1(n21331), .B0(n21215), .Y(n21616) );
  OAI21XL U24300 ( .A0(n6179), .A1(n21331), .B0(n21216), .Y(n21604) );
  OAI21XL U24301 ( .A0(n21223), .A1(n21222), .B0(n21221), .Y(n21230) );
  OAI21XL U24302 ( .A0(n21228), .A1(n21227), .B0(n21226), .Y(n21229) );
  INVX1 U24303 ( .A(n21862), .Y(n21266) );
  OAI21XL U24304 ( .A0(n6184), .A1(n21256), .B0(n21236), .Y(n21456) );
  NOR2X1 U24305 ( .A(n21266), .B(n21456), .Y(n21269) );
  OAI21XL U24306 ( .A0(n6213), .A1(n21256), .B0(n21238), .Y(n21475) );
  NOR2X1 U24307 ( .A(n21269), .B(n21239), .Y(n21272) );
  OAI21XL U24308 ( .A0(n25888), .A1(n21329), .B0(n21242), .Y(n21470) );
  OAI21XL U24309 ( .A0(n26140), .A1(n25887), .B0(w1[9]), .Y(n21244) );
  INVX1 U24310 ( .A(n21901), .Y(n21279) );
  OAI21XL U24311 ( .A0(n6207), .A1(n21311), .B0(n21248), .Y(n21513) );
  NOR2X1 U24312 ( .A(n21279), .B(n21513), .Y(n21282) );
  INVX1 U24313 ( .A(n21880), .Y(n21278) );
  OAI21XL U24314 ( .A0(n6209), .A1(n21256), .B0(n21250), .Y(n21461) );
  NOR2X1 U24315 ( .A(n21282), .B(n21251), .Y(n21285) );
  INVX1 U24316 ( .A(n21870), .Y(n21273) );
  OAI21XL U24317 ( .A0(n6183), .A1(n21256), .B0(n21253), .Y(n21457) );
  INVX1 U24318 ( .A(n21875), .Y(n21274) );
  OAI21XL U24319 ( .A0(n6211), .A1(n21256), .B0(n21255), .Y(n21460) );
  NOR2X1 U24320 ( .A(n21274), .B(n21460), .Y(n21277) );
  NAND2X1 U24321 ( .A(n21285), .B(n21258), .Y(n21287) );
  NOR2X1 U24322 ( .A(n21259), .B(n21287), .Y(n21290) );
  OAI21XL U24323 ( .A0(n21264), .A1(n21263), .B0(n21262), .Y(n21271) );
  OAI21XL U24324 ( .A0(n21269), .A1(n21268), .B0(n21267), .Y(n21270) );
  OAI21XL U24325 ( .A0(n21277), .A1(n21276), .B0(n21275), .Y(n21284) );
  OAI21XL U24326 ( .A0(n21282), .A1(n21281), .B0(n21280), .Y(n21283) );
  INVX1 U24327 ( .A(n21987), .Y(n21343) );
  OAI21XL U24328 ( .A0(n6166), .A1(n21311), .B0(n21293), .Y(n21508) );
  NOR2X1 U24329 ( .A(n21343), .B(n21508), .Y(n21346) );
  OAI21XL U24330 ( .A0(n26170), .A1(n21311), .B0(n21294), .Y(n21982) );
  INVX1 U24331 ( .A(n21982), .Y(n21342) );
  OAI21XL U24332 ( .A0(n6205), .A1(n21311), .B0(n21295), .Y(n21520) );
  NOR2X1 U24333 ( .A(n21346), .B(n21296), .Y(n21349) );
  OAI21XL U24334 ( .A0(n26172), .A1(n21311), .B0(n21297), .Y(n21961) );
  INVX1 U24335 ( .A(n21961), .Y(n21337) );
  OAI21XL U24336 ( .A0(n6187), .A1(n21311), .B0(n21298), .Y(n21514) );
  CLKINVX3 U24337 ( .A(n4631), .Y(n21333) );
  OAI21XL U24338 ( .A0(n6186), .A1(n21311), .B0(n21300), .Y(n21517) );
  OAI21XL U24339 ( .A0(n26160), .A1(n21333), .B0(n21303), .Y(n21426) );
  INVX1 U24340 ( .A(n21426), .Y(n21356) );
  OAI21X1 U24341 ( .A0(n6172), .A1(n21256), .B0(n21304), .Y(n21425) );
  NOR2X1 U24342 ( .A(n21356), .B(n21425), .Y(n21359) );
  OAI21XL U24343 ( .A0(n26166), .A1(n21333), .B0(n21305), .Y(n21422) );
  INVX1 U24344 ( .A(n21422), .Y(n21355) );
  NOR2X1 U24345 ( .A(n21359), .B(n21307), .Y(n21362) );
  OAI21XL U24346 ( .A0(n26167), .A1(n21311), .B0(n21308), .Y(n21992) );
  INVX1 U24347 ( .A(n21992), .Y(n21350) );
  OAI21XL U24348 ( .A0(n6215), .A1(n21311), .B0(n21309), .Y(n21509) );
  INVX1 U24349 ( .A(n21997), .Y(n21351) );
  OAI21XL U24350 ( .A0(n26141), .A1(n21333), .B0(n21312), .Y(n21511) );
  NOR2X1 U24351 ( .A(n21351), .B(n21511), .Y(n21354) );
  NAND2X1 U24352 ( .A(n21362), .B(n21314), .Y(n21364) );
  NOR2X1 U24353 ( .A(n21315), .B(n21364), .Y(n21336) );
  INVX1 U24354 ( .A(n21410), .Y(n21372) );
  NOR2X1 U24355 ( .A(n21372), .B(n21409), .Y(n21375) );
  INVX1 U24356 ( .A(n21406), .Y(n21371) );
  NOR2X1 U24357 ( .A(n21375), .B(n21320), .Y(n21378) );
  OAI21XL U24358 ( .A0(n26162), .A1(n21256), .B0(n21321), .Y(n21431) );
  INVX1 U24359 ( .A(n21431), .Y(n21366) );
  INVX1 U24360 ( .A(n21435), .Y(n21367) );
  NOR2X1 U24361 ( .A(n21367), .B(n21434), .Y(n21370) );
  NAND2X1 U24362 ( .A(n21378), .B(n21326), .Y(n21335) );
  INVX1 U24363 ( .A(n21418), .Y(n21380) );
  OR2X2 U24364 ( .A(n21380), .B(n21417), .Y(n21383) );
  OR2X2 U24365 ( .A(n21379), .B(n21413), .Y(n21334) );
  OAI21XL U24366 ( .A0(n21341), .A1(n21340), .B0(n21339), .Y(n21348) );
  OAI21XL U24367 ( .A0(n21346), .A1(n21345), .B0(n21344), .Y(n21347) );
  OAI21XL U24368 ( .A0(n21354), .A1(n21353), .B0(n21352), .Y(n21361) );
  OAI21XL U24369 ( .A0(n21359), .A1(n21358), .B0(n21357), .Y(n21360) );
  AOI21XL U24370 ( .A0(n21362), .A1(n21361), .B0(n21360), .Y(n21363) );
  OAI21XL U24371 ( .A0(n21370), .A1(n21369), .B0(n21368), .Y(n21377) );
  OAI21XL U24372 ( .A0(n21375), .A1(n21374), .B0(n21373), .Y(n21376) );
  AOI21XL U24373 ( .A0(n21378), .A1(n21377), .B0(n21376), .Y(n21386) );
  AOI21X1 U24374 ( .A0(n21383), .A1(n21382), .B0(n21381), .Y(n21384) );
  INVX4 U24375 ( .A(n21393), .Y(n21429) );
  INVX4 U24376 ( .A(n21429), .Y(n21628) );
  OAI21X2 U24377 ( .A0(n21628), .A1(n21379), .B0(n21394), .Y(n23413) );
  OAI21X2 U24378 ( .A0(n21628), .A1(n21372), .B0(n21395), .Y(n23394) );
  OAI21X2 U24379 ( .A0(n21628), .A1(n21371), .B0(n21396), .Y(n23230) );
  OAI21X2 U24380 ( .A0(n21519), .A1(n21367), .B0(n21397), .Y(n23406) );
  NAND2X1 U24381 ( .A(n3020), .B(n21430), .Y(n21398) );
  NAND2X1 U24382 ( .A(n21519), .B(n21425), .Y(n21399) );
  NAND2X1 U24383 ( .A(n23116), .B(n21421), .Y(n21400) );
  CMPR22X1 U24384 ( .A(n23394), .B(n21401), .CO(n22169), .S(n23393) );
  CMPR22X1 U24385 ( .A(n23230), .B(n21402), .CO(n21401), .S(n23229) );
  NAND2X1 U24386 ( .A(n21420), .B(n21380), .Y(n23398) );
  OAI21XL U24387 ( .A0(n21519), .A1(n21420), .B0(n21419), .Y(n23118) );
  MXI2X1 U24388 ( .A(y20[31]), .B(w1[31]), .S0(n21329), .Y(n23117) );
  NAND2X1 U24389 ( .A(n23420), .B(n21444), .Y(n21451) );
  CLKINVX3 U24390 ( .A(n21507), .Y(n21689) );
  CLKINVX3 U24391 ( .A(n21429), .Y(n23116) );
  OAI21XL U24392 ( .A0(n21689), .A1(n21731), .B0(n21459), .Y(n21561) );
  OAI21XL U24393 ( .A0(n21519), .A1(n21881), .B0(n21462), .Y(n21718) );
  OAI21XL U24394 ( .A0(n21689), .A1(n21698), .B0(n21463), .Y(n21570) );
  OAI21XL U24395 ( .A0(n21580), .A1(n21561), .B0(n21465), .Y(n21794) );
  OAI21XL U24396 ( .A0(n21689), .A1(n21683), .B0(n21472), .Y(n21558) );
  INVX1 U24397 ( .A(n21689), .Y(n21582) );
  NAND2XL U24398 ( .A(n23116), .B(n21844), .Y(n21474) );
  OAI21XL U24399 ( .A0(n21628), .A1(n21845), .B0(n21474), .Y(n21674) );
  CLKINVX3 U24400 ( .A(n21507), .Y(n21643) );
  NAND2XL U24401 ( .A(n23116), .B(n21852), .Y(n21476) );
  OAI21XL U24402 ( .A0(n21519), .A1(n21853), .B0(n21476), .Y(n21717) );
  AOI22XL U24403 ( .A0(n21582), .A1(n21674), .B0(n21643), .B1(n21717), .Y(
        n21563) );
  OAI21XL U24404 ( .A0(n21580), .A1(n21558), .B0(n21477), .Y(n21796) );
  OAI22XL U24405 ( .A0(n21794), .A1(n3172), .B0(n3096), .B1(n21796), .Y(n21633) );
  OAI21XL U24406 ( .A0(n21505), .A1(n21501), .B0(n21502), .Y(n21490) );
  OAI21XL U24407 ( .A0(n3020), .A1(n21993), .B0(n21510), .Y(n21711) );
  AOI22XL U24408 ( .A0(n21582), .A1(n21544), .B0(n21689), .B1(n21711), .Y(
        n21564) );
  OAI21XL U24409 ( .A0(n3020), .A1(n21998), .B0(n21512), .Y(n21709) );
  OAI21XL U24410 ( .A0(n21519), .A1(n21962), .B0(n21515), .Y(n21671) );
  OAI21XL U24411 ( .A0(n21689), .A1(n21728), .B0(n21516), .Y(n21567) );
  OAI21XL U24412 ( .A0(n21519), .A1(n21978), .B0(n21518), .Y(n21708) );
  OAI21XL U24413 ( .A0(n3020), .A1(n21983), .B0(n21521), .Y(n21678) );
  OAI21XL U24414 ( .A0(n21689), .A1(n21523), .B0(n21522), .Y(n21566) );
  OAI21XL U24415 ( .A0(n21580), .A1(n21567), .B0(n21525), .Y(n21795) );
  OAI21XL U24416 ( .A0(n21689), .A1(n21714), .B0(n21533), .Y(n21585) );
  AOI22XL U24417 ( .A0(n21507), .A1(n21718), .B0(n21643), .B1(n21534), .Y(
        n21591) );
  NAND2XL U24418 ( .A(n21580), .B(n21591), .Y(n21535) );
  OAI21XL U24419 ( .A0(n21580), .A1(n21585), .B0(n21535), .Y(n21602) );
  OAI21XL U24420 ( .A0(n21689), .A1(n21699), .B0(n21536), .Y(n21583) );
  OAI21XL U24421 ( .A0(n21689), .A1(n21539), .B0(n21538), .Y(n21588) );
  OAI21XL U24422 ( .A0(n21580), .A1(n21583), .B0(n21541), .Y(n21607) );
  OAI22XL U24423 ( .A0(n21602), .A1(n3172), .B0(n3096), .B1(n21607), .Y(n21650) );
  AOI22XL U24424 ( .A0(n21507), .A1(n21711), .B0(n21643), .B1(n21709), .Y(
        n21592) );
  OAI21XL U24425 ( .A0(n21689), .A1(n21543), .B0(n21542), .Y(n21589) );
  OAI21XL U24426 ( .A0(n21689), .A1(n21546), .B0(n21545), .Y(n21594) );
  OAI21XL U24427 ( .A0(n21580), .A1(n21589), .B0(n21548), .Y(n21603) );
  NAND2XL U24428 ( .A(n3020), .B(n21578), .Y(n21555) );
  NAND2XL U24429 ( .A(n21519), .B(n21600), .Y(n21557) );
  OAI21XL U24430 ( .A0(n21628), .A1(n21601), .B0(n21557), .Y(n21684) );
  AOI22XL U24431 ( .A0(n21507), .A1(n21697), .B0(n21643), .B1(n21684), .Y(
        n21629) );
  AOI22XL U24432 ( .A0(n3095), .A1(n21629), .B0(n21559), .B1(n21580), .Y(
        n21763) );
  AOI22XL U24433 ( .A0(n21763), .A1(n3172), .B0(n21767), .B1(n3096), .Y(n21665) );
  AOI21XL U24434 ( .A0(n21665), .A1(n3037), .B0(n21803), .Y(n21574) );
  OAI21XL U24435 ( .A0(n21580), .A1(n21566), .B0(n21565), .Y(n21768) );
  OAI21XL U24436 ( .A0(n21580), .A1(n21570), .B0(n21569), .Y(n21766) );
  AOI22XL U24437 ( .A0(n21582), .A1(n21684), .B0(n21643), .B1(n21581), .Y(
        n21606) );
  AOI22XL U24438 ( .A0(n3095), .A1(n21606), .B0(n21584), .B1(n21580), .Y(
        n21777) );
  OAI21XL U24439 ( .A0(n21580), .A1(n21588), .B0(n21587), .Y(n21780) );
  AOI21XL U24440 ( .A0(n21751), .A1(n3037), .B0(n21803), .Y(n21596) );
  OAI21XL U24441 ( .A0(n21580), .A1(n21594), .B0(n21593), .Y(n21782) );
  OAI22XL U24442 ( .A0(n21603), .A1(n21560), .B0(n3096), .B1(n21602), .Y(
        n21867) );
  NAND2XL U24443 ( .A(n3020), .B(n21616), .Y(n21605) );
  OAI21XL U24444 ( .A0(n21628), .A1(n21617), .B0(n21605), .Y(n21721) );
  AOI22XL U24445 ( .A0(n3095), .A1(n21745), .B0(n21606), .B1(n21580), .Y(
        n21646) );
  OAI21XL U24446 ( .A0(n21867), .A1(n3037), .B0(n21610), .Y(n21611) );
  INVXL U24447 ( .A(n21700), .Y(n21622) );
  INVXL U24448 ( .A(n21701), .Y(n21621) );
  AOI22XL U24449 ( .A0(n21582), .A1(n21622), .B0(n21643), .B1(n21621), .Y(
        n21660) );
  NAND2XL U24450 ( .A(n21519), .B(n21775), .Y(n21624) );
  OAI21XL U24451 ( .A0(n21628), .A1(n21776), .B0(n21624), .Y(n21719) );
  AOI22XL U24452 ( .A0(n21582), .A1(n21719), .B0(n21643), .B1(n21644), .Y(
        n21662) );
  AOI22XL U24453 ( .A0(n3095), .A1(n21660), .B0(n21662), .B1(n21580), .Y(
        n21630) );
  NAND2XL U24454 ( .A(n21519), .B(n21809), .Y(n21627) );
  OAI21XL U24455 ( .A0(n21628), .A1(n21810), .B0(n21627), .Y(n21688) );
  AOI22XL U24456 ( .A0(n21507), .A1(n21688), .B0(n21643), .B1(n21721), .Y(
        n21661) );
  AOI22XL U24457 ( .A0(n21630), .A1(n3172), .B0(n21798), .B1(n3096), .Y(n21631) );
  AOI21XL U24458 ( .A0(n21631), .A1(n3037), .B0(n21803), .Y(n21632) );
  OAI21XL U24459 ( .A0(n3037), .A1(n21633), .B0(n21632), .Y(n21634) );
  OAI21XL U24460 ( .A0(n21635), .A1(n21801), .B0(n21634), .Y(n21636) );
  OR2X2 U24461 ( .A(n21757), .B(n21756), .Y(n22127) );
  NAND2XL U24462 ( .A(n21643), .B(n21719), .Y(n21642) );
  OAI21XL U24463 ( .A0(n21689), .A1(n21701), .B0(n21642), .Y(n21743) );
  AOI22XL U24464 ( .A0(n21507), .A1(n21644), .B0(n21643), .B1(n21688), .Y(
        n21746) );
  AOI22XL U24465 ( .A0(n3095), .A1(n21645), .B0(n21746), .B1(n21580), .Y(
        n21647) );
  AOI22XL U24466 ( .A0(n21647), .A1(n21560), .B0(n21646), .B1(n3096), .Y(
        n21648) );
  AOI21XL U24467 ( .A0(n21648), .A1(n3037), .B0(n21803), .Y(n21649) );
  OAI21XL U24468 ( .A0(n3037), .A1(n21650), .B0(n21649), .Y(n21651) );
  OAI21XL U24469 ( .A0(n21652), .A1(n21801), .B0(n21651), .Y(n21653) );
  AOI21XL U24470 ( .A0(n21655), .A1(n3222), .B0(n21849), .Y(n21654) );
  AOI22XL U24471 ( .A0(n21663), .A1(n3172), .B0(n21764), .B1(n3096), .Y(n21664) );
  AOI21XL U24472 ( .A0(n21664), .A1(n3037), .B0(n21803), .Y(n21667) );
  NAND2XL U24473 ( .A(n21665), .B(n3171), .Y(n21666) );
  OAI21XL U24474 ( .A0(n21668), .A1(n21787), .B0(n3222), .Y(n21670) );
  AOI211XL U24475 ( .A0(n21672), .A1(n21671), .B0(n21697), .C0(n21719), .Y(
        n21682) );
  NAND2XL U24476 ( .A(n3095), .B(n21507), .Y(n21696) );
  OAI21XL U24477 ( .A0(n3037), .A1(n21707), .B0(n21801), .Y(n21675) );
  AOI21XL U24478 ( .A0(n21675), .A1(n21674), .B0(n21673), .Y(n21681) );
  AOI21XL U24479 ( .A0(n3037), .A1(n21582), .B0(n21676), .Y(n21679) );
  AOI211XL U24480 ( .A0(n3037), .A1(n3095), .B0(n21793), .C0(n21801), .Y(
        n21677) );
  OAI21XL U24481 ( .A0(n21679), .A1(n21678), .B0(n21677), .Y(n21680) );
  NOR2XL U24482 ( .A(n21803), .B(n3096), .Y(n21687) );
  AOI211XL U24483 ( .A0(n21687), .A1(n3095), .B0(n21686), .C0(n21702), .Y(
        n21694) );
  OAI21XL U24484 ( .A0(n21722), .A1(n21689), .B0(n21688), .Y(n21692) );
  NAND2XL U24485 ( .A(n3096), .B(n21580), .Y(n21690) );
  AOI22XL U24486 ( .A0(n21692), .A1(n21691), .B0(n21702), .B1(n21690), .Y(
        n21693) );
  AOI22XL U24487 ( .A0(n21710), .A1(n21697), .B0(n21744), .B1(n21580), .Y(
        n21706) );
  AOI211XL U24488 ( .A0(n21793), .A1(n21783), .B0(n21698), .C0(n21801), .Y(
        n21705) );
  NAND2XL U24489 ( .A(n3171), .B(n3096), .Y(n21716) );
  AOI21XL U24490 ( .A0(n21716), .A1(n21801), .B0(n21699), .Y(n21704) );
  AOI22XL U24491 ( .A0(n21702), .A1(n3172), .B0(n21701), .B1(n21700), .Y(
        n21703) );
  AOI22XL U24492 ( .A0(n21710), .A1(n21709), .B0(n21720), .B1(n21708), .Y(
        n21715) );
  OAI21XL U24493 ( .A0(n21712), .A1(n21711), .B0(n3171), .Y(n21713) );
  AOI31XL U24494 ( .A0(n21715), .A1(n21714), .A2(n21713), .B0(n21801), .Y(
        n21726) );
  AOI21XL U24495 ( .A0(n21793), .A1(n3095), .B0(n21801), .Y(n21727) );
  OAI21XL U24496 ( .A0(n21716), .A1(n3095), .B0(n21801), .Y(n21730) );
  AOI22XL U24497 ( .A0(n21722), .A1(n21721), .B0(n21720), .B1(n21719), .Y(
        n21724) );
  NAND4BXL U24498 ( .AN(n21726), .B(n21725), .C(n21724), .D(n21723), .Y(n21735) );
  AOI211XL U24499 ( .A0(n21793), .A1(n21507), .B0(n21729), .C0(n21728), .Y(
        n21734) );
  AOI211XL U24500 ( .A0(n21801), .A1(n21582), .B0(n21732), .C0(n21731), .Y(
        n21733) );
  INVXL U24501 ( .A(n22195), .Y(n21740) );
  AOI22XL U24502 ( .A0(n3095), .A1(n21744), .B0(n21580), .B1(n21743), .Y(
        n21748) );
  OAI21XL U24503 ( .A0(n3096), .A1(n21748), .B0(n21747), .Y(n21749) );
  OAI21XL U24504 ( .A0(n21749), .A1(n3171), .B0(n21801), .Y(n21750) );
  AOI21XL U24505 ( .A0(n3171), .A1(n21751), .B0(n21750), .Y(n21752) );
  AOI21XL U24506 ( .A0(n21877), .A1(n21803), .B0(n21752), .Y(n21753) );
  OAI21XL U24507 ( .A0(n21854), .A1(n21755), .B0(n21754), .Y(n22130) );
  AOI22XL U24508 ( .A0(n21764), .A1(n3172), .B0(n21763), .B1(n3096), .Y(n21765) );
  AOI21XL U24509 ( .A0(n21765), .A1(n3037), .B0(n21803), .Y(n21771) );
  AOI21XL U24510 ( .A0(n21774), .A1(n3222), .B0(n21849), .Y(n21773) );
  AOI22XL U24511 ( .A0(n21778), .A1(n21560), .B0(n21777), .B1(n3096), .Y(
        n21779) );
  AOI21XL U24512 ( .A0(n21779), .A1(n3037), .B0(n21803), .Y(n21785) );
  AOI21XL U24513 ( .A0(n21789), .A1(n3222), .B0(n21849), .Y(n21788) );
  OAI22XL U24514 ( .A0(n21795), .A1(n21560), .B0(n3096), .B1(n21794), .Y(
        n21858) );
  AOI22XL U24515 ( .A0(n21798), .A1(n3172), .B0(n21797), .B1(n3096), .Y(n21799) );
  OAI21XL U24516 ( .A0(n21858), .A1(n3037), .B0(n21800), .Y(n21802) );
  AOI22XL U24517 ( .A0(n21804), .A1(n21803), .B0(n21802), .B1(n21801), .Y(
        n21806) );
  OAI21XL U24518 ( .A0(n21952), .A1(n22107), .B0(n21953), .Y(n21835) );
  OAI21XL U24519 ( .A0(n21856), .A1(n3096), .B0(n3171), .Y(n21857) );
  OAI21XL U24520 ( .A0(n21865), .A1(n3096), .B0(n3171), .Y(n21866) );
  OAI21XL U24521 ( .A0(n21925), .A1(n21934), .B0(n21926), .Y(n21890) );
  OAI21XL U24522 ( .A0(n21912), .A1(n21917), .B0(n21913), .Y(n22042) );
  AOI21XL U24523 ( .A0(n22048), .A1(n22039), .B0(n22042), .Y(n21896) );
  OAI21XL U24524 ( .A0(n22051), .A1(n21897), .B0(n21896), .Y(n21907) );
  NOR2X1 U24525 ( .A(n21904), .B(n21903), .Y(n22044) );
  OAI21XL U24526 ( .A0(n22051), .A1(n21911), .B0(n21910), .Y(n21916) );
  OAI21XL U24527 ( .A0(n22051), .A1(n21963), .B0(n21970), .Y(n21920) );
  AOI21XL U24528 ( .A0(n21931), .A1(n21935), .B0(n21922), .Y(n21923) );
  OAI21XL U24529 ( .A0(n22051), .A1(n21924), .B0(n21923), .Y(n21929) );
  OAI21XL U24530 ( .A0(n22051), .A1(n21933), .B0(n21932), .Y(n21937) );
  OAI21XL U24531 ( .A0(n22051), .A1(n21943), .B0(n21944), .Y(n21942) );
  OAI21XL U24532 ( .A0(n21949), .A1(n22106), .B0(n22107), .Y(n21950) );
  OAI21XL U24533 ( .A0(n22052), .A1(n22043), .B0(n22053), .Y(n21966) );
  OR2X2 U24534 ( .A(n22058), .B(n22018), .Y(n22022) );
  OAI21XL U24535 ( .A0(n22071), .A1(n22064), .B0(n22072), .Y(n22007) );
  OAI21XL U24536 ( .A0(n22057), .A1(n22018), .B0(n22014), .Y(n22015) );
  OAI21XL U24537 ( .A0(n22070), .A1(n22026), .B0(n22025), .Y(n22029) );
  OAI21XL U24538 ( .A0(n22070), .A1(n22035), .B0(n22036), .Y(n22034) );
  OAI21XL U24539 ( .A0(n22045), .A1(n22044), .B0(n22043), .Y(n22046) );
  OAI21XL U24540 ( .A0(n22051), .A1(n22050), .B0(n22049), .Y(n22056) );
  OAI21XL U24541 ( .A0(n22070), .A1(n22058), .B0(n22057), .Y(n22062) );
  AOI21XL U24542 ( .A0(n22067), .A1(n22066), .B0(n22065), .Y(n22068) );
  OAI21XL U24543 ( .A0(n22070), .A1(n22069), .B0(n22068), .Y(n22075) );
  CMPR22X1 U24544 ( .A(n23406), .B(n22076), .CO(n21402), .S(n23405) );
  OAI21XL U24545 ( .A0(n22092), .A1(n22079), .B0(n22078), .Y(n22084) );
  OAI21XL U24546 ( .A0(n22092), .A1(n22085), .B0(n22089), .Y(n22088) );
  XNOR2X1 U24547 ( .A(n22088), .B(n22087), .Y(n22302) );
  AOI21XL U24548 ( .A0(n22128), .A1(n22127), .B0(n22094), .Y(n22097) );
  XOR2X1 U24549 ( .A(n22097), .B(n22096), .Y(n22202) );
  AOI21XL U24550 ( .A0(n22117), .A1(n22102), .B0(n22098), .Y(n22101) );
  AOI21XL U24551 ( .A0(n22117), .A1(n22105), .B0(n22104), .Y(n22110) );
  OAI21XL U24552 ( .A0(n22114), .A1(n22113), .B0(n22112), .Y(n22115) );
  AOI21XL U24553 ( .A0(n22117), .A1(n22116), .B0(n22115), .Y(n22120) );
  CMPR22X1 U24554 ( .A(n23402), .B(n22125), .CO(n22076), .S(n23401) );
  XNOR2XL U24555 ( .A(n22132), .B(n22131), .Y(n22185) );
  OAI21XL U24556 ( .A0(n22135), .A1(n22134), .B0(n22133), .Y(n22137) );
  AOI2BB1X2 U24557 ( .A0N(n22149), .A1N(n22254), .B0(n22333), .Y(n22150) );
  AOI2BB1X2 U24558 ( .A0N(n22150), .A1N(n22252), .B0(n22421), .Y(n22151) );
  AOI2BB1X2 U24559 ( .A0N(n22151), .A1N(n22256), .B0(n22448), .Y(n22152) );
  OAI21XL U24560 ( .A0(n22203), .A1(n22185), .B0(n22153), .Y(n22154) );
  OAI21XL U24561 ( .A0(n22158), .A1(n22157), .B0(n22156), .Y(n22159) );
  CMPR22X1 U24562 ( .A(n23420), .B(n23409), .CO(n22125), .S(n23417) );
  CMPR22X1 U24563 ( .A(n23413), .B(n22169), .CO(n22170), .S(n23412) );
  CMPR22X1 U24564 ( .A(n23398), .B(n22170), .CO(n22171), .S(n23397) );
  CMPR32X1 U24565 ( .A(n23405), .B(n3082), .C(n22177), .CO(n22180), .S(n23404)
         );
  ADDFHX1 U24566 ( .A(n23401), .B(n3079), .CI(n22178), .CO(n22177), .S(n23400)
         );
  CMPR32X1 U24567 ( .A(n22179), .B(n22395), .C(n23417), .CO(n22178), .S(n23416) );
  ADDFHX1 U24568 ( .A(n23229), .B(n22461), .CI(n22180), .CO(n22176), .S(n22181) );
  NAND4BXL U24569 ( .AN(n22201), .B(n22252), .C(n22421), .D(n22256), .Y(n22211) );
  INVXL U24570 ( .A(n23420), .Y(n22221) );
  INVXL U24571 ( .A(n23230), .Y(n22220) );
  INVXL U24572 ( .A(n23402), .Y(n22219) );
  INVXL U24573 ( .A(n23394), .Y(n22218) );
  NAND4XL U24574 ( .A(n22221), .B(n22220), .C(n22219), .D(n22218), .Y(n22226)
         );
  NOR2XL U24575 ( .A(n23413), .B(n23406), .Y(n22224) );
  INVXL U24576 ( .A(n23398), .Y(n22223) );
  NAND3XL U24577 ( .A(n22224), .B(n22223), .C(n22222), .Y(n22225) );
  NOR2X1 U24578 ( .A(n22226), .B(n22225), .Y(n23129) );
  OAI21XL U24579 ( .A0(n3126), .A1(n22232), .B0(n22231), .Y(n22318) );
  OAI21XL U24580 ( .A0(n3126), .A1(n22234), .B0(n22233), .Y(n22317) );
  OAI21XL U24581 ( .A0(n3126), .A1(n22236), .B0(n22235), .Y(n22316) );
  OAI21XL U24582 ( .A0(n22343), .A1(n22316), .B0(n22238), .Y(n22406) );
  OAI21XL U24583 ( .A0(n3126), .A1(n22241), .B0(n22240), .Y(n22322) );
  OAI21XL U24584 ( .A0(n3126), .A1(n22243), .B0(n22242), .Y(n22326) );
  OAI22XL U24585 ( .A0(n22426), .A1(n22322), .B0(n22326), .B1(n3129), .Y(
        n22413) );
  NOR2XL U24586 ( .A(n3126), .B(n22277), .Y(n22245) );
  AOI21XL U24587 ( .A0(n22292), .A1(n3126), .B0(n22245), .Y(n22320) );
  NOR2XL U24588 ( .A(n3126), .B(n22246), .Y(n22249) );
  AOI22XL U24589 ( .A0(n22320), .A1(n22343), .B0(n22324), .B1(n3129), .Y(
        n22368) );
  OAI21XL U24590 ( .A0(n3130), .A1(n22413), .B0(n22251), .Y(n22266) );
  NOR2XL U24591 ( .A(n22266), .B(n3082), .Y(n22265) );
  OAI21XL U24592 ( .A0(n3126), .A1(n22423), .B0(n22253), .Y(n22437) );
  OAI21XL U24593 ( .A0(n3126), .A1(n22335), .B0(n22255), .Y(n22323) );
  OAI22XL U24594 ( .A0(n22343), .A1(n22437), .B0(n22323), .B1(n3129), .Y(
        n22411) );
  OAI21XL U24595 ( .A0(n3126), .A1(n22450), .B0(n22257), .Y(n22436) );
  NAND2XL U24596 ( .A(n3126), .B(n22448), .Y(n22259) );
  OAI21XL U24597 ( .A0(n22261), .A1(n6168), .B0(n3082), .Y(n22262) );
  NOR2XL U24598 ( .A(n22267), .B(n3082), .Y(n22269) );
  OAI21XL U24599 ( .A0(n3126), .A1(n22275), .B0(n22274), .Y(n22331) );
  NOR2XL U24600 ( .A(n3126), .B(n22276), .Y(n22279) );
  NAND2XL U24601 ( .A(n22342), .B(n22426), .Y(n22280) );
  OAI21XL U24602 ( .A0(n22426), .A1(n22331), .B0(n22280), .Y(n22375) );
  NOR2XL U24603 ( .A(n3126), .B(n22283), .Y(n22284) );
  AOI21XL U24604 ( .A0(n22285), .A1(n3126), .B0(n22284), .Y(n22338) );
  OAI21XL U24605 ( .A0(n3126), .A1(n22289), .B0(n22288), .Y(n22332) );
  NOR2XL U24606 ( .A(n22332), .B(n3129), .Y(n22290) );
  OAI21XL U24607 ( .A0(n3079), .A1(n22375), .B0(n22291), .Y(n22313) );
  NOR2XL U24608 ( .A(n3126), .B(n22293), .Y(n22294) );
  OAI21XL U24609 ( .A0(n3126), .A1(n22299), .B0(n22298), .Y(n22341) );
  OAI21XL U24610 ( .A0(n3126), .A1(n22304), .B0(n22303), .Y(n22340) );
  NAND2XL U24611 ( .A(n22397), .B(n22426), .Y(n22311) );
  OAI21XL U24612 ( .A0(n22250), .A1(n22340), .B0(n22311), .Y(n22372) );
  OAI21XL U24613 ( .A0(n22315), .A1(n22461), .B0(n22314), .Y(n23311) );
  AOI21XL U24614 ( .A0(n22320), .A1(n22395), .B0(n22319), .Y(n22362) );
  OAI21XL U24615 ( .A0(n22361), .A1(n3079), .B0(n22321), .Y(n22390) );
  NOR2XL U24616 ( .A(n22390), .B(n3082), .Y(n22330) );
  OAI22XL U24617 ( .A0(n22426), .A1(n22323), .B0(n22322), .B1(n3129), .Y(
        n22440) );
  OAI21XL U24618 ( .A0(n22440), .A1(n3130), .B0(n3082), .Y(n22328) );
  OAI21XL U24619 ( .A0(n22343), .A1(n22326), .B0(n22325), .Y(n22364) );
  NOR2XL U24620 ( .A(n22364), .B(n3079), .Y(n22327) );
  AOI22XL U24621 ( .A0(n22396), .A1(n22426), .B0(n22397), .B1(n3129), .Y(
        n22354) );
  OAI22XL U24622 ( .A0(n22426), .A1(n22332), .B0(n22331), .B1(n3129), .Y(
        n22353) );
  NOR2XL U24623 ( .A(n3126), .B(n22334), .Y(n22337) );
  AOI22XL U24624 ( .A0(n22338), .A1(n22426), .B0(n22427), .B1(n22395), .Y(
        n22455) );
  AOI21XL U24625 ( .A0(n22455), .A1(n3079), .B0(n22124), .Y(n22339) );
  OAI21XL U24626 ( .A0(n3079), .A1(n22353), .B0(n22339), .Y(n22347) );
  OAI22XL U24627 ( .A0(n22426), .A1(n22341), .B0(n22340), .B1(n3129), .Y(
        n22356) );
  OAI21XL U24628 ( .A0(n22356), .A1(n3079), .B0(n22345), .Y(n22385) );
  OAI21XL U24629 ( .A0(n22418), .A1(n22349), .B0(n22348), .Y(n23305) );
  OAI21XL U24630 ( .A0(n3130), .A1(n22353), .B0(n22352), .Y(n22447) );
  OAI21XL U24631 ( .A0(n3130), .A1(n22356), .B0(n22355), .Y(n22392) );
  NOR2XL U24632 ( .A(n22392), .B(n3082), .Y(n22357) );
  OAI21XL U24633 ( .A0(n3130), .A1(n22361), .B0(n22360), .Y(n22393) );
  NAND2XL U24634 ( .A(n22362), .B(n3130), .Y(n22363) );
  OAI21XL U24635 ( .A0(n3130), .A1(n22364), .B0(n22363), .Y(n22444) );
  OAI21XL U24636 ( .A0(n22372), .A1(n3130), .B0(n22371), .Y(n22394) );
  NOR2XL U24637 ( .A(n22394), .B(n3082), .Y(n22377) );
  OAI21XL U24638 ( .A0(n3130), .A1(n22375), .B0(n22374), .Y(n22433) );
  NAND2XL U24639 ( .A(n22381), .B(n22124), .Y(n22382) );
  NOR2XL U24640 ( .A(n22386), .B(n3082), .Y(n22387) );
  NOR2XL U24641 ( .A(n22397), .B(n22426), .Y(n22400) );
  NAND2XL U24642 ( .A(n22402), .B(n3130), .Y(n22404) );
  NOR2X1 U24643 ( .A(n22409), .B(n23244), .Y(n23383) );
  OAI21XL U24644 ( .A0(n3079), .A1(n22413), .B0(n22412), .Y(n22416) );
  NAND2XL U24645 ( .A(n22414), .B(n22124), .Y(n22415) );
  AOI21XL U24646 ( .A0(n22454), .A1(n3129), .B0(n3130), .Y(n22429) );
  AOI21XL U24647 ( .A0(n22429), .A1(n22428), .B0(n22124), .Y(n22430) );
  OAI21XL U24648 ( .A0(n22433), .A1(n3082), .B0(n22432), .Y(n22434) );
  OAI21XL U24649 ( .A0(n22435), .A1(n22461), .B0(n22434), .Y(n23380) );
  OAI21XL U24650 ( .A0(n22439), .A1(n22438), .B0(n3082), .Y(n22442) );
  OAI21XL U24651 ( .A0(n22444), .A1(n3082), .B0(n22443), .Y(n22445) );
  OAI21XL U24652 ( .A0(n22446), .A1(n22461), .B0(n22445), .Y(n23374) );
  INVXL U24653 ( .A(n22458), .Y(n22459) );
  AOI21XL U24654 ( .A0(n23044), .A1(n3216), .B0(n22469), .Y(n2099) );
  NOR2XL U24655 ( .A(n26311), .B(n23063), .Y(n23062) );
  NAND2XL U24656 ( .A(iter[2]), .B(n23062), .Y(n23055) );
  NOR2XL U24657 ( .A(n26309), .B(n23055), .Y(n23054) );
  NAND2XL U24658 ( .A(iter[4]), .B(n23054), .Y(n23058) );
  NOR2XL U24659 ( .A(n26312), .B(n23058), .Y(n23057) );
  NAND2XL U24660 ( .A(iter[6]), .B(n23057), .Y(n23060) );
  OAI21XL U24661 ( .A0(learning_rate[23]), .A1(n25856), .B0(n24007), .Y(n22470) );
  OAI21XL U24662 ( .A0(n22472), .A1(n26195), .B0(n25230), .Y(n22473) );
  AOI21XL U24663 ( .A0(n3223), .A1(sigma10[31]), .B0(n22473), .Y(n22475) );
  OAI21XL U24664 ( .A0(n4583), .A1(n26313), .B0(n25236), .Y(n22474) );
  NAND2XL U24665 ( .A(n3111), .B(data[95]), .Y(n22480) );
  CMPR32X1 U24666 ( .A(n22490), .B(n22621), .C(n10775), .CO(M6_mult_x_15_n545), 
        .S(M6_mult_x_15_n546) );
  AND3X2 U24667 ( .A(n22512), .B(n22511), .C(n22493), .Y(n22891) );
  OAI21XL U24668 ( .A0(n11082), .A1(n22894), .B0(n22494), .Y(n22495) );
  OAI21XL U24669 ( .A0(n22506), .A1(n22499), .B0(n22498), .Y(n22529) );
  OAI21XL U24670 ( .A0(n22800), .A1(n22909), .B0(n22502), .Y(n22503) );
  OAI21XL U24671 ( .A0(n22506), .A1(n22505), .B0(n22504), .Y(n22516) );
  OAI21XL U24672 ( .A0(n23091), .A1(n22909), .B0(n22509), .Y(n22510) );
  NOR2X4 U24673 ( .A(n22512), .B(n22511), .Y(n22892) );
  OAI21XL U24674 ( .A0(n22800), .A1(n22894), .B0(n22513), .Y(n22514) );
  OAI21XL U24675 ( .A0(n23095), .A1(n22909), .B0(n22520), .Y(n22521) );
  OAI21XL U24676 ( .A0(n22913), .A1(n22894), .B0(n22522), .Y(n22523) );
  OAI21XL U24677 ( .A0(n23091), .A1(n22894), .B0(n22524), .Y(n22525) );
  OAI21XL U24678 ( .A0(n23098), .A1(n22894), .B0(n22535), .Y(n22536) );
  OAI21XL U24679 ( .A0(n23095), .A1(n22894), .B0(n22537), .Y(n22538) );
  OAI21XL U24680 ( .A0(n22913), .A1(n22984), .B0(n22539), .Y(n22540) );
  OAI21XL U24681 ( .A0(n11082), .A1(n22909), .B0(n22541), .Y(n22542) );
  CMPR32X1 U24682 ( .A(n22549), .B(M6_mult_x_15_n464), .C(n22543), .CO(
        M6_mult_x_15_n458), .S(M6_mult_x_15_n459) );
  OAI21XL U24683 ( .A0(n23098), .A1(n22909), .B0(n22544), .Y(n22545) );
  OAI21XL U24684 ( .A0(n22800), .A1(n11089), .B0(n22546), .Y(n22547) );
  CMPR32X1 U24685 ( .A(n11063), .B(n22549), .C(n22548), .CO(M6_mult_x_15_n452), 
        .S(M6_mult_x_15_n453) );
  OAI21XL U24686 ( .A0(n23076), .A1(n22894), .B0(n22551), .Y(n22552) );
  OAI21XL U24687 ( .A0(n23101), .A1(n22894), .B0(n22560), .Y(n22561) );
  NOR2X4 U24688 ( .A(n22563), .B(n22562), .Y(n22988) );
  OAI21XL U24689 ( .A0(n23076), .A1(n22984), .B0(n22565), .Y(n22566) );
  OAI21XL U24690 ( .A0(n23104), .A1(n22894), .B0(n22571), .Y(n22572) );
  OAI21XL U24691 ( .A0(n23095), .A1(n22984), .B0(n22573), .Y(n22574) );
  OAI21XL U24692 ( .A0(n22643), .A1(n22582), .B0(n22584), .Y(n22775) );
  OAI21XL U24693 ( .A0(n23026), .A1(n23154), .B0(n22577), .Y(n22578) );
  CMPR32X1 U24694 ( .A(n11058), .B(n22636), .C(n22579), .CO(M6_mult_x_15_n495), 
        .S(M6_mult_x_15_n496) );
  OAI21XL U24695 ( .A0(n11082), .A1(n23025), .B0(n22580), .Y(n22581) );
  OAI21XL U24696 ( .A0(n22643), .A1(n22589), .B0(n22588), .Y(n22632) );
  OAI21XL U24697 ( .A0(n23107), .A1(n22894), .B0(n22597), .Y(n22598) );
  OAI21XL U24698 ( .A0(n22913), .A1(n23005), .B0(n22599), .Y(n22600) );
  OAI21XL U24699 ( .A0(n22643), .A1(n22604), .B0(n22603), .Y(n22762) );
  CLKINVX3 U24700 ( .A(n22896), .Y(n22953) );
  AOI222XL U24701 ( .A0(n22953), .A1(n11059), .B0(n10797), .B1(n11058), .C0(
        n22952), .C1(n23151), .Y(n22607) );
  OAI21XL U24702 ( .A0(n23139), .A1(n22834), .B0(n22607), .Y(n22608) );
  AOI222XL U24703 ( .A0(n23023), .A1(n10775), .B0(n22887), .B1(n10769), .C0(
        n23021), .C1(n23002), .Y(n22609) );
  OAI21XL U24704 ( .A0(n22993), .A1(n23025), .B0(n22609), .Y(n22610) );
  XOR2XL U24705 ( .A(n22610), .B(n3054), .Y(M6_mult_x_15_n1157) );
  OAI21XL U24706 ( .A0(n23139), .A1(n23005), .B0(n22611), .Y(n22612) );
  OAI21XL U24707 ( .A0(n23095), .A1(n23025), .B0(n22613), .Y(n22615) );
  OAI21XL U24708 ( .A0(n23098), .A1(n23005), .B0(n22616), .Y(n22617) );
  AOI222XL U24709 ( .A0(n22953), .A1(n23151), .B0(n10797), .B1(n10789), .C0(
        n22952), .C1(n3220), .Y(n22618) );
  OAI21XL U24710 ( .A0(n23155), .A1(n22834), .B0(n22618), .Y(n22619) );
  XOR2XL U24711 ( .A(n22619), .B(n3221), .Y(M6_mult_x_15_n1207) );
  OAI21XL U24712 ( .A0(n23095), .A1(n22834), .B0(n22620), .Y(n22622) );
  OAI21XL U24713 ( .A0(n23091), .A1(n22834), .B0(n22623), .Y(n22624) );
  OAI21XL U24714 ( .A0(n23095), .A1(n22912), .B0(n22625), .Y(n22626) );
  OAI21XL U24715 ( .A0(n23104), .A1(n22909), .B0(n22627), .Y(n22628) );
  OAI21XL U24716 ( .A0(n23111), .A1(n22894), .B0(n22633), .Y(n22634) );
  CMPR32X1 U24717 ( .A(n22636), .B(M6_mult_x_15_n513), .C(n22635), .CO(
        M6_mult_x_15_n504), .S(M6_mult_x_15_n505) );
  AOI222XL U24718 ( .A0(n22932), .A1(n10789), .B0(n22904), .B1(n3220), .C0(
        n22931), .C1(n26496), .Y(n22637) );
  OAI21XL U24719 ( .A0(n23148), .A1(n22912), .B0(n22637), .Y(n22638) );
  XOR2XL U24720 ( .A(n22638), .B(n3053), .Y(M6_mult_x_15_n1181) );
  OAI21XL U24721 ( .A0(n23098), .A1(n23025), .B0(n22639), .Y(n22640) );
  OAI21XL U24722 ( .A0(n22643), .A1(n22642), .B0(n22641), .Y(n22648) );
  AOI222XL U24723 ( .A0(n22953), .A1(n11058), .B0(n10797), .B1(n23151), .C0(
        n22952), .C1(n10789), .Y(n22649) );
  OAI21XL U24724 ( .A0(n23142), .A1(n22834), .B0(n22649), .Y(n22650) );
  XOR2XL U24725 ( .A(n22650), .B(n3221), .Y(M6_mult_x_15_n1206) );
  AOI222XL U24726 ( .A0(n22932), .A1(n26496), .B0(n22904), .B1(n10775), .C0(
        n22931), .C1(n10769), .Y(n22651) );
  OAI21XL U24727 ( .A0(n22924), .A1(n22912), .B0(n22651), .Y(n22652) );
  XOR2XL U24728 ( .A(n22652), .B(n3053), .Y(M6_mult_x_15_n1183) );
  OAI21XL U24729 ( .A0(n23104), .A1(n22984), .B0(n22653), .Y(n22654) );
  OAI21XL U24730 ( .A0(n11082), .A1(n23005), .B0(n22655), .Y(n22656) );
  AOI222XL U24731 ( .A0(n23023), .A1(n26496), .B0(n22887), .B1(n10775), .C0(
        n23021), .C1(n10769), .Y(n22657) );
  OAI21XL U24732 ( .A0(n22924), .A1(n23025), .B0(n22657), .Y(n22658) );
  XOR2XL U24733 ( .A(n22658), .B(n3054), .Y(M6_mult_x_15_n1156) );
  AOI222XL U24734 ( .A0(n23023), .A1(n10769), .B0(n22887), .B1(n23002), .C0(
        n23021), .C1(n10749), .Y(n22659) );
  OAI21XL U24735 ( .A0(n22998), .A1(n23025), .B0(n22659), .Y(n22660) );
  XOR2XL U24736 ( .A(n22660), .B(n3054), .Y(M6_mult_x_15_n1158) );
  AOI222XL U24737 ( .A0(n23023), .A1(n11058), .B0(n22887), .B1(n23151), .C0(
        n23021), .C1(n10789), .Y(n22661) );
  OAI21XL U24738 ( .A0(n23142), .A1(n23025), .B0(n22661), .Y(n22662) );
  XOR2XL U24739 ( .A(n22662), .B(n3054), .Y(M6_mult_x_15_n1152) );
  AOI222XL U24740 ( .A0(n22932), .A1(n23151), .B0(n22904), .B1(n10789), .C0(
        n22931), .C1(n3220), .Y(n22663) );
  OAI21XL U24741 ( .A0(n23155), .A1(n22912), .B0(n22663), .Y(n22664) );
  XOR2XL U24742 ( .A(n22664), .B(n3053), .Y(M6_mult_x_15_n1180) );
  AOI222XL U24743 ( .A0(n22953), .A1(n3219), .B0(n10797), .B1(n11073), .C0(
        n22952), .C1(n11063), .Y(n22665) );
  OAI21XL U24744 ( .A0(n23101), .A1(n22834), .B0(n22665), .Y(n22666) );
  OAI21XL U24745 ( .A0(n23026), .A1(n22894), .B0(n22667), .Y(n22668) );
  OAI21XL U24746 ( .A0(n22800), .A1(n23005), .B0(n22669), .Y(n22670) );
  AOI222XL U24747 ( .A0(n23023), .A1(n3220), .B0(n22887), .B1(n22867), .C0(
        n23021), .C1(n10775), .Y(n22671) );
  OAI21XL U24748 ( .A0(n22869), .A1(n23025), .B0(n22671), .Y(n22672) );
  XOR2XL U24749 ( .A(n22672), .B(n3054), .Y(M6_mult_x_15_n1155) );
  AOI222XL U24750 ( .A0(n22932), .A1(n3220), .B0(n22904), .B1(n22867), .C0(
        n22931), .C1(n10775), .Y(n22673) );
  OAI21XL U24751 ( .A0(n22869), .A1(n22912), .B0(n22673), .Y(n22674) );
  XOR2XL U24752 ( .A(n22674), .B(n3053), .Y(M6_mult_x_15_n1182) );
  OAI21XL U24753 ( .A0(n22800), .A1(n22984), .B0(n22675), .Y(n22676) );
  OAI21XL U24754 ( .A0(n23142), .A1(n22984), .B0(n22677), .Y(n22678) );
  AOI222XL U24755 ( .A0(n23023), .A1(n11059), .B0(n22887), .B1(n11058), .C0(
        n23021), .C1(n23151), .Y(n22679) );
  OAI21XL U24756 ( .A0(n23139), .A1(n23025), .B0(n22679), .Y(n22680) );
  XOR2XL U24757 ( .A(n22680), .B(n3054), .Y(M6_mult_x_15_n1151) );
  OAI21XL U24758 ( .A0(n11082), .A1(n22834), .B0(n22681), .Y(n22682) );
  AOI222XL U24759 ( .A0(n23023), .A1(n23002), .B0(n22887), .B1(n10749), .C0(
        n23021), .C1(n3116), .Y(n22683) );
  OAI21XL U24760 ( .A0(n23006), .A1(n23025), .B0(n22683), .Y(n22684) );
  XOR2XL U24761 ( .A(n22684), .B(n3054), .Y(M6_mult_x_15_n1159) );
  OAI21XL U24762 ( .A0(n23091), .A1(n23005), .B0(n22685), .Y(n22686) );
  OAI21XL U24763 ( .A0(n23098), .A1(n22834), .B0(n22687), .Y(n22688) );
  AOI222XL U24764 ( .A0(n22932), .A1(n11058), .B0(n22904), .B1(n23151), .C0(
        n22931), .C1(n10789), .Y(n22689) );
  OAI21XL U24765 ( .A0(n23142), .A1(n22912), .B0(n22689), .Y(n22690) );
  OAI21XL U24766 ( .A0(n23139), .A1(n22984), .B0(n22691), .Y(n22692) );
  AOI222XL U24767 ( .A0(n22953), .A1(n11073), .B0(n10797), .B1(n11063), .C0(
        n22952), .C1(n23109), .Y(n22693) );
  OAI21XL U24768 ( .A0(n23104), .A1(n22834), .B0(n22693), .Y(n22694) );
  XOR2XL U24769 ( .A(n22694), .B(n3221), .Y(M6_mult_x_15_n1199) );
  OAI21XL U24770 ( .A0(n23107), .A1(n22912), .B0(n22695), .Y(n22696) );
  OAI21XL U24771 ( .A0(n22978), .A1(n22909), .B0(n22697), .Y(n22699) );
  OAI21XL U24772 ( .A0(n22985), .A1(n22909), .B0(n22703), .Y(n22704) );
  OAI21XL U24773 ( .A0(n22909), .A1(n22989), .B0(n4706), .Y(n22705) );
  OAI21XL U24774 ( .A0(n22978), .A1(n22894), .B0(n22706), .Y(n22707) );
  OAI21XL U24775 ( .A0(n22985), .A1(n22894), .B0(n22711), .Y(n22712) );
  OAI21XL U24776 ( .A0(n22894), .A1(n22989), .B0(n4708), .Y(n22714) );
  OAI21XL U24777 ( .A0(n22993), .A1(n22909), .B0(n22715), .Y(n22717) );
  CMPR22X1 U24778 ( .A(n22719), .B(n22718), .CO(n23046), .S(n23032) );
  OAI21XL U24779 ( .A0(n22998), .A1(n22909), .B0(n22720), .Y(n22721) );
  CMPR22X1 U24780 ( .A(n3119), .B(n22722), .CO(n22718), .S(n23035) );
  OAI21XL U24781 ( .A0(n23006), .A1(n22909), .B0(n22723), .Y(n22724) );
  CMPR22X1 U24782 ( .A(n22726), .B(n22725), .CO(n23033), .S(M6_mult_x_15_n672)
         );
  CMPR32X1 U24783 ( .A(n22729), .B(n22728), .C(n22727), .CO(M6_mult_x_15_n641), 
        .S(M6_mult_x_15_n642) );
  OAI21XL U24784 ( .A0(n23091), .A1(n22912), .B0(n22730), .Y(n22731) );
  OAI21XL U24785 ( .A0(n22993), .A1(n22894), .B0(n22732), .Y(n22733) );
  OAI21XL U24786 ( .A0(n23091), .A1(n23025), .B0(n22734), .Y(n22735) );
  OAI21XL U24787 ( .A0(n23155), .A1(n22984), .B0(n22736), .Y(n22738) );
  AOI222XL U24788 ( .A0(n23023), .A1(n10789), .B0(n22887), .B1(n3220), .C0(
        n23021), .C1(n26496), .Y(n22739) );
  OAI21XL U24789 ( .A0(n23148), .A1(n23025), .B0(n22739), .Y(n22740) );
  XOR2XL U24790 ( .A(n22740), .B(n3054), .Y(M6_mult_x_15_n1154) );
  OAI21XL U24791 ( .A0(n22869), .A1(n22909), .B0(n22741), .Y(n22742) );
  OAI21XL U24792 ( .A0(n22993), .A1(n22984), .B0(n22743), .Y(n22744) );
  OAI21XL U24793 ( .A0(n23091), .A1(n22984), .B0(n22745), .Y(n22746) );
  OAI21XL U24794 ( .A0(n23095), .A1(n23005), .B0(n22747), .Y(n22748) );
  OAI21XL U24795 ( .A0(n23098), .A1(n22984), .B0(n22749), .Y(n22750) );
  AOI222XL U24796 ( .A0(n23023), .A1(n23151), .B0(n22887), .B1(n10789), .C0(
        n23021), .C1(n3220), .Y(n22751) );
  OAI21XL U24797 ( .A0(n23155), .A1(n23025), .B0(n22751), .Y(n22752) );
  OAI21XL U24798 ( .A0(n23111), .A1(n22909), .B0(n22753), .Y(n22754) );
  OAI21XL U24799 ( .A0(n23148), .A1(n22894), .B0(n22755), .Y(n22756) );
  OAI21XL U24800 ( .A0(n22869), .A1(n22894), .B0(n22757), .Y(n22758) );
  AOI222XL U24801 ( .A0(n23023), .A1(n26493), .B0(n22887), .B1(n11059), .C0(
        n23021), .C1(n11058), .Y(n22768) );
  OAI21XL U24802 ( .A0(n23145), .A1(n23025), .B0(n22768), .Y(n22769) );
  OAI21XL U24803 ( .A0(n22800), .A1(n22912), .B0(n22770), .Y(n22771) );
  AOI222XL U24804 ( .A0(n22932), .A1(n11062), .B0(n22904), .B1(n3217), .C0(
        n22931), .C1(n26493), .Y(n22781) );
  OAI21XL U24805 ( .A0(n23135), .A1(n22912), .B0(n22781), .Y(n22782) );
  OAI21XL U24806 ( .A0(n11082), .A1(n22912), .B0(n22783), .Y(n22784) );
  OAI21XL U24807 ( .A0(n23101), .A1(n22984), .B0(n22785), .Y(n22786) );
  OAI21XL U24808 ( .A0(n23142), .A1(n22909), .B0(n22787), .Y(n22788) );
  OAI21XL U24809 ( .A0(n22800), .A1(n23025), .B0(n22789), .Y(n22790) );
  OAI21XL U24810 ( .A0(n23139), .A1(n22909), .B0(n22791), .Y(n22792) );
  OAI21XL U24811 ( .A0(n23101), .A1(n22909), .B0(n22793), .Y(n22794) );
  AOI222XL U24812 ( .A0(n22953), .A1(n3217), .B0(n10797), .B1(n23022), .C0(
        n22952), .C1(n11059), .Y(n22795) );
  OAI21XL U24813 ( .A0(n23026), .A1(n22834), .B0(n22795), .Y(n22796) );
  AOI222XL U24814 ( .A0(n22953), .A1(n26493), .B0(n10797), .B1(n11059), .C0(
        n22952), .C1(n11058), .Y(n22797) );
  OAI21XL U24815 ( .A0(n23145), .A1(n22834), .B0(n22797), .Y(n22798) );
  OAI21XL U24816 ( .A0(n22800), .A1(n22834), .B0(n22799), .Y(n22801) );
  OAI21XL U24817 ( .A0(n23104), .A1(n23005), .B0(n22802), .Y(n22803) );
  OAI21XL U24818 ( .A0(n23026), .A1(n23005), .B0(n22804), .Y(n22805) );
  AOI222XL U24819 ( .A0(n22953), .A1(n23109), .B0(n10797), .B1(n11062), .C0(
        n22952), .C1(n3217), .Y(n22806) );
  OAI21XL U24820 ( .A0(n23111), .A1(n22834), .B0(n22806), .Y(n22807) );
  OAI21XL U24821 ( .A0(n23148), .A1(n22984), .B0(n22808), .Y(n22809) );
  OAI21XL U24822 ( .A0(n23098), .A1(n22912), .B0(n22810), .Y(n22811) );
  OAI21XL U24823 ( .A0(n23135), .A1(n22894), .B0(n22812), .Y(n22813) );
  AOI222XL U24824 ( .A0(n22932), .A1(n11059), .B0(n22904), .B1(n11058), .C0(
        n22931), .C1(n23151), .Y(n22814) );
  OAI21XL U24825 ( .A0(n23139), .A1(n22912), .B0(n22814), .Y(n22815) );
  OAI21XL U24826 ( .A0(n23148), .A1(n22909), .B0(n22816), .Y(n22817) );
  OAI21XL U24827 ( .A0(n23104), .A1(n23025), .B0(n22818), .Y(n22819) );
  AOI222XL U24828 ( .A0(n22953), .A1(n11063), .B0(n10797), .B1(n23109), .C0(
        n22952), .C1(n11062), .Y(n22820) );
  OAI21XL U24829 ( .A0(n23107), .A1(n22834), .B0(n22820), .Y(n22821) );
  AOI222XL U24830 ( .A0(n23003), .A1(n10789), .B0(n22969), .B1(n3220), .C0(
        n23001), .C1(n26496), .Y(n22822) );
  OAI21XL U24831 ( .A0(n23148), .A1(n23005), .B0(n22822), .Y(n22823) );
  XOR2XL U24832 ( .A(n22823), .B(n3055), .Y(M6_mult_x_15_n1127) );
  OAI21XL U24833 ( .A0(n23107), .A1(n22909), .B0(n22824), .Y(n22825) );
  OAI21XL U24834 ( .A0(n22993), .A1(n23154), .B0(n22826), .Y(n22827) );
  CMPR32X1 U24835 ( .A(n10749), .B(n3221), .C(n22828), .CO(M6_mult_x_15_n578), 
        .S(M6_mult_x_15_n579) );
  OAI21XL U24836 ( .A0(n22913), .A1(n23025), .B0(n22829), .Y(n22830) );
  OAI21XL U24837 ( .A0(n23145), .A1(n22894), .B0(n22831), .Y(n22832) );
  OAI21XL U24838 ( .A0(n22913), .A1(n22834), .B0(n22833), .Y(n22835) );
  OAI21XL U24839 ( .A0(n23107), .A1(n23005), .B0(n22836), .Y(n22837) );
  OAI21XL U24840 ( .A0(n23076), .A1(n23005), .B0(n22839), .Y(n22840) );
  OAI21XL U24841 ( .A0(n23026), .A1(n22984), .B0(n22841), .Y(n22842) );
  AOI222XL U24842 ( .A0(n23003), .A1(n3220), .B0(n22969), .B1(n22867), .C0(
        n23001), .C1(n10775), .Y(n22843) );
  OAI21XL U24843 ( .A0(n22869), .A1(n23005), .B0(n22843), .Y(n22844) );
  XOR2XL U24844 ( .A(n22844), .B(n3055), .Y(M6_mult_x_15_n1128) );
  AOI222XL U24845 ( .A0(n22932), .A1(n3217), .B0(n22904), .B1(n23022), .C0(
        n22931), .C1(n11059), .Y(n22845) );
  OAI21XL U24846 ( .A0(n23026), .A1(n22912), .B0(n22845), .Y(n22846) );
  XOR2XL U24847 ( .A(n22846), .B(n3053), .Y(M6_mult_x_15_n1176) );
  OAI21XL U24848 ( .A0(n22869), .A1(n22984), .B0(n22847), .Y(n22848) );
  OAI21XL U24849 ( .A0(n23111), .A1(n22984), .B0(n22849), .Y(n22850) );
  OAI21XL U24850 ( .A0(n23101), .A1(n23025), .B0(n22851), .Y(n22852) );
  OAI21XL U24851 ( .A0(n23135), .A1(n22909), .B0(n22853), .Y(n22854) );
  OAI21XL U24852 ( .A0(n23145), .A1(n22984), .B0(n22855), .Y(n22856) );
  OAI21XL U24853 ( .A0(n22998), .A1(n22894), .B0(n22857), .Y(n22858) );
  OAI21XL U24854 ( .A0(n23111), .A1(n23025), .B0(n22859), .Y(n22860) );
  OAI21XL U24855 ( .A0(n23135), .A1(n22984), .B0(n22861), .Y(n22862) );
  OAI21XL U24856 ( .A0(n23107), .A1(n23025), .B0(n22863), .Y(n22864) );
  OAI21XL U24857 ( .A0(n23135), .A1(n23005), .B0(n22865), .Y(n22866) );
  OAI21XL U24858 ( .A0(n22869), .A1(n23154), .B0(n22868), .Y(n22870) );
  CMPR32X1 U24859 ( .A(n3221), .B(n10769), .C(n22871), .CO(M6_mult_x_15_n556), 
        .S(M6_mult_x_15_n557) );
  OAI21XL U24860 ( .A0(n23104), .A1(n22912), .B0(n22872), .Y(n22873) );
  OAI21XL U24861 ( .A0(n23155), .A1(n22894), .B0(n22874), .Y(n22875) );
  OAI21XL U24862 ( .A0(n22924), .A1(n22894), .B0(n22876), .Y(n22877) );
  OAI21XL U24863 ( .A0(n23155), .A1(n22909), .B0(n22878), .Y(n22879) );
  AOI222XL U24864 ( .A0(n22932), .A1(n26493), .B0(n22904), .B1(n11059), .C0(
        n22931), .C1(n11058), .Y(n22880) );
  OAI21XL U24865 ( .A0(n23145), .A1(n22912), .B0(n22880), .Y(n22881) );
  OAI21XL U24866 ( .A0(n23142), .A1(n22894), .B0(n22882), .Y(n22883) );
  OAI21XL U24867 ( .A0(n23139), .A1(n22894), .B0(n22884), .Y(n22885) );
  OAI21XL U24868 ( .A0(n23076), .A1(n23025), .B0(n22889), .Y(n22890) );
  OAI21XL U24869 ( .A0(n23006), .A1(n22894), .B0(n22893), .Y(n22895) );
  OAI21XL U24870 ( .A0(n23076), .A1(n22834), .B0(n22899), .Y(n22900) );
  OAI21XL U24871 ( .A0(n23101), .A1(n22912), .B0(n22901), .Y(n22902) );
  OAI21XL U24872 ( .A0(n23076), .A1(n22912), .B0(n22906), .Y(n22907) );
  OAI21XL U24873 ( .A0(n23026), .A1(n22909), .B0(n22908), .Y(n22910) );
  OAI21XL U24874 ( .A0(n22913), .A1(n22912), .B0(n22911), .Y(n22914) );
  OAI21XL U24875 ( .A0(n22998), .A1(n22984), .B0(n22915), .Y(n22916) );
  AOI222XL U24876 ( .A0(n22988), .A1(n23002), .B0(n22980), .B1(n10749), .C0(
        n22976), .C1(n3116), .Y(n22917) );
  OAI21XL U24877 ( .A0(n23006), .A1(n22984), .B0(n22917), .Y(n22918) );
  OAI21XL U24878 ( .A0(n23101), .A1(n23005), .B0(n22919), .Y(n22920) );
  OAI21XL U24879 ( .A0(n22924), .A1(n22984), .B0(n22921), .Y(n22922) );
  OAI21XL U24880 ( .A0(n22924), .A1(n23154), .B0(n22923), .Y(n22925) );
  CMPR32X1 U24881 ( .A(n3221), .B(n23002), .C(n22926), .CO(M6_mult_x_15_n567), 
        .S(M6_mult_x_15_n568) );
  OAI21XL U24882 ( .A0(n23145), .A1(n22909), .B0(n22929), .Y(n22930) );
  OAI21XL U24883 ( .A0(n23111), .A1(n22912), .B0(n22933), .Y(n22934) );
  AOI222XL U24884 ( .A0(n22988), .A1(n11063), .B0(n22980), .B1(n23109), .C0(
        n22976), .C1(n11062), .Y(n22935) );
  OAI21XL U24885 ( .A0(n23107), .A1(n22984), .B0(n22935), .Y(n22936) );
  OAI21XL U24886 ( .A0(n23142), .A1(n23005), .B0(n22937), .Y(n22938) );
  OAI21XL U24887 ( .A0(n22978), .A1(n23154), .B0(n22939), .Y(n22940) );
  OAI21XL U24888 ( .A0(n22985), .A1(n23154), .B0(n22942), .Y(n22943) );
  OAI21XL U24889 ( .A0(n22998), .A1(n23154), .B0(n22944), .Y(n22945) );
  OAI21XL U24890 ( .A0(n23006), .A1(n23154), .B0(n22946), .Y(n22947) );
  CMPR22X1 U24891 ( .A(n22949), .B(n22948), .CO(n22958), .S(M6_mult_x_15_n612)
         );
  CMPR32X1 U24892 ( .A(n3116), .B(n22951), .C(n22950), .CO(M6_mult_x_15_n589), 
        .S(M6_mult_x_15_n590) );
  AOI222XL U24893 ( .A0(n22953), .A1(n11062), .B0(n10797), .B1(n3217), .C0(
        n22952), .C1(n26493), .Y(n22954) );
  OAI21XL U24894 ( .A0(n23135), .A1(n22834), .B0(n22954), .Y(n22955) );
  OAI21XL U24895 ( .A0(n23135), .A1(n23025), .B0(n22956), .Y(n22957) );
  CMPR32X1 U24896 ( .A(n22987), .B(n22959), .C(n22958), .CO(n22950), .S(
        M6_mult_x_15_n601) );
  CMPR22X1 U24897 ( .A(n22961), .B(n22960), .CO(n22948), .S(M6_mult_x_15_n623)
         );
  OAI21XL U24898 ( .A0(n23145), .A1(n23005), .B0(n22962), .Y(n22963) );
  OAI21XL U24899 ( .A0(n23111), .A1(n23005), .B0(n22964), .Y(n22965) );
  AOI222XL U24900 ( .A0(n23003), .A1(n10749), .B0(n22969), .B1(n3116), .C0(
        n23001), .C1(n22987), .Y(n22966) );
  OAI21XL U24901 ( .A0(n22978), .A1(n23005), .B0(n22966), .Y(n22968) );
  INVXL U24902 ( .A(n22971), .Y(n22972) );
  OAI21XL U24903 ( .A0(n22985), .A1(n23005), .B0(n22972), .Y(n22973) );
  OAI21XL U24904 ( .A0(n23005), .A1(n22989), .B0(n22974), .Y(n22975) );
  OAI21XL U24905 ( .A0(n22978), .A1(n22984), .B0(n22977), .Y(n22979) );
  INVXL U24906 ( .A(n22982), .Y(n22983) );
  OAI21XL U24907 ( .A0(n22985), .A1(n22984), .B0(n22983), .Y(n22986) );
  OAI21XL U24908 ( .A0(n22984), .A1(n22989), .B0(n4705), .Y(n22991) );
  AOI222XL U24909 ( .A0(n23003), .A1(n10775), .B0(n22969), .B1(n10769), .C0(
        n23001), .C1(n23002), .Y(n22992) );
  OAI21XL U24910 ( .A0(n22993), .A1(n23005), .B0(n22992), .Y(n22994) );
  XOR2XL U24911 ( .A(n22994), .B(n3055), .Y(n23011) );
  CMPR22X1 U24912 ( .A(n22996), .B(n22995), .CO(n23028), .S(n23015) );
  AOI222XL U24913 ( .A0(n23003), .A1(n10769), .B0(n22969), .B1(n23002), .C0(
        n23001), .C1(n10749), .Y(n22997) );
  OAI21XL U24914 ( .A0(n22998), .A1(n23005), .B0(n22997), .Y(n22999) );
  XOR2XL U24915 ( .A(n22999), .B(n3055), .Y(n23014) );
  CMPR22X1 U24916 ( .A(n3056), .B(n23000), .CO(n22995), .S(n23018) );
  AOI222XL U24917 ( .A0(n23003), .A1(n23002), .B0(n22969), .B1(n10749), .C0(
        n23001), .C1(n3116), .Y(n23004) );
  OAI21XL U24918 ( .A0(n23006), .A1(n23005), .B0(n23004), .Y(n23007) );
  CMPR22X1 U24919 ( .A(n23009), .B(n23008), .CO(n23016), .S(M6_mult_x_15_n714)
         );
  CMPR32X1 U24920 ( .A(n23012), .B(n23011), .C(n23010), .CO(M6_mult_x_15_n692), 
        .S(M6_mult_x_15_n693) );
  CMPR32X1 U24921 ( .A(n23015), .B(n23014), .C(n23013), .CO(n23010), .S(
        M6_mult_x_15_n700) );
  CMPR32X1 U24922 ( .A(n23018), .B(n23017), .C(n23016), .CO(n23013), .S(
        M6_mult_x_15_n707) );
  CMPR22X1 U24923 ( .A(n23020), .B(n23019), .CO(n23008), .S(M6_mult_x_15_n719)
         );
  OAI21XL U24924 ( .A0(n23026), .A1(n23025), .B0(n23024), .Y(n23027) );
  CMPR22X1 U24925 ( .A(n23029), .B(n23028), .CO(M6_mult_x_15_n694), .S(n23012)
         );
  CMPR32X1 U24926 ( .A(n23032), .B(n23031), .C(n23030), .CO(n22727), .S(
        M6_mult_x_15_n652) );
  CMPR32X1 U24927 ( .A(n23035), .B(n23034), .C(n23033), .CO(n23030), .S(
        M6_mult_x_15_n662) );
  CMPR22X1 U24928 ( .A(n23037), .B(n23036), .CO(n22725), .S(M6_mult_x_15_n680)
         );
  AND2XL U24929 ( .A(M2_U3_U1_enc_tree_1__1__12_), .B(
        M2_U3_U1_enc_tree_1__1__14_), .Y(n25984) );
  AND2XL U24930 ( .A(M2_U4_U1_enc_tree_1__1__12_), .B(
        M2_U4_U1_enc_tree_1__1__14_), .Y(n25989) );
  NOR2XL U24931 ( .A(n21256), .B(cs[2]), .Y(n23071) );
  AOI21XL U24932 ( .A0(n23038), .A1(n23235), .B0(n23133), .Y(n23043) );
  CMPR22X1 U24933 ( .A(n3055), .B(n23045), .CO(n23019), .S(M6_mult_x_15_n724)
         );
  CMPR22X1 U24934 ( .A(n23047), .B(n23046), .CO(M6_mult_x_15_n643), .S(n22729)
         );
  CMPR22X1 U24935 ( .A(n3058), .B(n23048), .CO(n23036), .S(M6_mult_x_15_n688)
         );
  NAND2XL U24936 ( .A(y20[11]), .B(n2972), .Y(n2512) );
  NAND2XL U24937 ( .A(y20[22]), .B(n2972), .Y(n2501) );
  NAND2XL U24938 ( .A(y20[8]), .B(n2972), .Y(n2515) );
  NAND2XL U24939 ( .A(y20[16]), .B(n2972), .Y(n2507) );
  NAND2XL U24940 ( .A(y20[23]), .B(n2972), .Y(n2500) );
  NAND2XL U24941 ( .A(y20[17]), .B(n2972), .Y(n2506) );
  NAND2XL U24942 ( .A(y20[15]), .B(n2972), .Y(n2508) );
  NAND2XL U24943 ( .A(y20[4]), .B(n2972), .Y(n2519) );
  NAND2XL U24944 ( .A(y20[5]), .B(n2972), .Y(n2518) );
  NAND2XL U24945 ( .A(y20[18]), .B(n2972), .Y(n2505) );
  NAND2XL U24946 ( .A(y20[14]), .B(n2972), .Y(n2509) );
  NAND2XL U24947 ( .A(y20[31]), .B(n2972), .Y(n2492) );
  NAND2XL U24948 ( .A(y20[12]), .B(n2972), .Y(n2511) );
  NAND2XL U24949 ( .A(y20[10]), .B(n2972), .Y(n2513) );
  NAND2XL U24950 ( .A(y20[7]), .B(n2972), .Y(n2516) );
  NAND2XL U24951 ( .A(y20[6]), .B(n2972), .Y(n2517) );
  NAND2XL U24952 ( .A(y20[19]), .B(n2972), .Y(n2504) );
  NAND2XL U24953 ( .A(y20[13]), .B(n2972), .Y(n2510) );
  NAND2XL U24954 ( .A(y20[21]), .B(n2972), .Y(n2502) );
  NAND2XL U24955 ( .A(y20[20]), .B(n2972), .Y(n2503) );
  NAND2XL U24956 ( .A(y20[30]), .B(n2972), .Y(n2493) );
  NAND2XL U24957 ( .A(y20[26]), .B(n2972), .Y(n2497) );
  NAND2XL U24958 ( .A(y20[29]), .B(n2972), .Y(n2494) );
  NAND2XL U24959 ( .A(y20[25]), .B(n2972), .Y(n2498) );
  NAND2XL U24960 ( .A(y20[24]), .B(n2972), .Y(n2499) );
  NAND2XL U24961 ( .A(y20[27]), .B(n2972), .Y(n2496) );
  NAND2XL U24962 ( .A(y20[28]), .B(n2972), .Y(n2495) );
  NAND2XL U24963 ( .A(n2972), .B(y20[3]), .Y(n2520) );
  NAND2XL U24964 ( .A(n2972), .B(y20[2]), .Y(n2521) );
  NAND2XL U24965 ( .A(n2972), .B(y20[0]), .Y(n2523) );
  NAND2XL U24966 ( .A(n2972), .B(y20[9]), .Y(n2514) );
  NAND2XL U24967 ( .A(n2972), .B(y20[1]), .Y(n2522) );
  NAND2XL U24968 ( .A(in_valid_d), .B(n25886), .Y(n23969) );
  INVXL U24969 ( .A(valid[1]), .Y(n23974) );
  OAI22XL U24970 ( .A0(n23969), .A1(n23049), .B0(n25664), .B1(n23974), .Y(N40)
         );
  NAND2XL U24971 ( .A(n24015), .B(n24008), .Y(n23052) );
  NAND2XL U24972 ( .A(n23051), .B(learning_rate[27]), .Y(n23050) );
  OAI21XL U24973 ( .A0(learning_rate[27]), .A1(n23051), .B0(n23050), .Y(n23982) );
  AOI21XL U24974 ( .A0(n26309), .A1(n23055), .B0(n23054), .Y(n23056) );
  NAND2XL U24975 ( .A(n23985), .B(n23056), .Y(n1744) );
  AOI21XL U24976 ( .A0(n26312), .A1(n23058), .B0(n23057), .Y(n23059) );
  NAND2XL U24977 ( .A(n23985), .B(n23059), .Y(n1746) );
  NOR2XL U24978 ( .A(n26308), .B(n23060), .Y(n25858) );
  AOI21XL U24979 ( .A0(n26308), .A1(n23060), .B0(n25858), .Y(n23061) );
  NAND2XL U24980 ( .A(n23985), .B(n23061), .Y(n1748) );
  AOI21XL U24981 ( .A0(n26311), .A1(n23063), .B0(n23062), .Y(n23064) );
  NAND2XL U24982 ( .A(n23985), .B(n23064), .Y(n1742) );
  INVXL U24983 ( .A(n24007), .Y(n23068) );
  NOR2XL U24984 ( .A(n23065), .B(n23980), .Y(n23066) );
  OAI21XL U24985 ( .A0(n23066), .A1(n24003), .B0(n24008), .Y(n23067) );
  AOI22XL U24986 ( .A0(n23068), .A1(n23067), .B0(n23980), .B1(n23985), .Y(
        n2627) );
  AOI211XL U24987 ( .A0(n25428), .A1(n7885), .B0(n23970), .C0(n25886), .Y(
        n23070) );
  NOR2XL U24988 ( .A(n23969), .B(cs[1]), .Y(n23069) );
  AOI211XL U24989 ( .A0(n3120), .A1(n23974), .B0(n23070), .C0(n23069), .Y(
        n2491) );
  OAI222XL U24990 ( .A0(n3117), .A1(w1[172]), .B0(n3226), .B1(w1[300]), .C0(
        w1[204]), .C1(n3228), .Y(n1928) );
  OAI222XL U24991 ( .A0(n3117), .A1(w1[32]), .B0(n3226), .B1(w1[160]), .C0(
        w1[64]), .C1(n3228), .Y(n1752) );
  OAI21XL U24992 ( .A0(n23076), .A1(n11089), .B0(n23075), .Y(n23077) );
  NAND2XL U24993 ( .A(n3111), .B(data[63]), .Y(n23080) );
  AOI22XL U24994 ( .A0(n21166), .A1(sigma10[31]), .B0(in_valid_t), .B1(w2[31]), 
        .Y(n23079) );
  OAI21XL U24995 ( .A0(n3045), .A1(n26310), .B0(n23085), .Y(n23086) );
  OAI21XL U24996 ( .A0(n23091), .A1(n11089), .B0(n23090), .Y(n23092) );
  OAI21XL U24997 ( .A0(n23095), .A1(n11089), .B0(n23094), .Y(n23096) );
  OAI21XL U24998 ( .A0(n23098), .A1(n11089), .B0(n23097), .Y(n23099) );
  OAI21XL U24999 ( .A0(n23101), .A1(n11089), .B0(n23100), .Y(n23102) );
  OAI21XL U25000 ( .A0(n23104), .A1(n11089), .B0(n23103), .Y(n23105) );
  OAI21XL U25001 ( .A0(n23107), .A1(n11089), .B0(n23106), .Y(n23108) );
  OAI21XL U25002 ( .A0(n23111), .A1(n11089), .B0(n23110), .Y(n23112) );
  AOI22XL U25003 ( .A0(n3042), .A1(n23117), .B0(n23116), .B1(n23115), .Y(
        n23131) );
  NAND4XL U25004 ( .A(n23121), .B(n23120), .C(n23119), .D(n23118), .Y(n23127)
         );
  NAND4XL U25005 ( .A(n23125), .B(n23124), .C(n23123), .D(n23122), .Y(n23126)
         );
  NOR2XL U25006 ( .A(n23127), .B(n23126), .Y(n23128) );
  OAI21XL U25007 ( .A0(n23129), .A1(n23128), .B0(n3222), .Y(n23130) );
  AOI222XL U25008 ( .A0(n23137), .A1(n23429), .B0(in_valid_t), .B1(target[31]), 
        .C0(n23428), .C1(target_temp[31]), .Y(n2263) );
  OAI21XL U25009 ( .A0(n23135), .A1(n11089), .B0(n23134), .Y(n23136) );
  OAI21XL U25010 ( .A0(n23139), .A1(n23154), .B0(n23138), .Y(n23140) );
  OAI21XL U25011 ( .A0(n23142), .A1(n23154), .B0(n23141), .Y(n23143) );
  OAI21XL U25012 ( .A0(n23145), .A1(n11089), .B0(n23144), .Y(n23146) );
  OAI21XL U25013 ( .A0(n23148), .A1(n23154), .B0(n23147), .Y(n23149) );
  OAI21XL U25014 ( .A0(n23155), .A1(n23154), .B0(n23153), .Y(n23156) );
  NAND4XL U25015 ( .A(n23160), .B(n23159), .C(n23158), .D(n23157), .Y(n23166)
         );
  NAND4XL U25016 ( .A(n23164), .B(n23163), .C(n23162), .D(n23161), .Y(n23165)
         );
  NOR2XL U25017 ( .A(n23166), .B(n23165), .Y(n23167) );
  AOI22XL U25018 ( .A0(n3101), .A1(n23170), .B0(n15008), .B1(n23169), .Y(
        n23171) );
  INVXL U25019 ( .A(M1_U4_U1_or2_tree_0__1__28_), .Y(M1_U4_U1_or2_inv_0__28_)
         );
  INVXL U25020 ( .A(M1_U4_U1_or2_tree_0__2__24_), .Y(M1_U4_U1_or2_inv_0__24_)
         );
  INVXL U25021 ( .A(M1_U4_U1_or2_tree_0__1__20_), .Y(M1_U4_U1_or2_inv_0__20_)
         );
  INVXL U25022 ( .A(M1_U3_U1_or2_tree_0__1__28_), .Y(M1_U3_U1_or2_inv_0__28_)
         );
  INVXL U25023 ( .A(M1_a_5_), .Y(M1_U3_U1_or2_inv_0__26_) );
  INVXL U25024 ( .A(M1_U3_U1_or2_tree_0__2__24_), .Y(M1_U3_U1_or2_inv_0__24_)
         );
  INVXL U25025 ( .A(n4567), .Y(M1_U3_U1_or2_inv_0__22_) );
  INVXL U25026 ( .A(M1_U3_U1_or2_tree_0__1__20_), .Y(M1_U3_U1_or2_inv_0__20_)
         );
  INVXL U25027 ( .A(M1_a_13_), .Y(M1_U3_U1_or2_inv_0__18_) );
  INVXL U25028 ( .A(M1_a_17_), .Y(M1_U3_U1_or2_inv_0__14_) );
  INVXL U25029 ( .A(M1_a_21_), .Y(M1_U3_U1_or2_inv_0__10_) );
  INVXL U25030 ( .A(M1_U4_U1_enc_tree_1__1__28_), .Y(M1_U4_U1_or2_inv_1__28_)
         );
  INVXL U25031 ( .A(M1_U4_U1_or2_tree_1__2__24_), .Y(M1_U4_U1_or2_inv_1__24_)
         );
  INVXL U25032 ( .A(M1_U4_U1_enc_tree_1__1__20_), .Y(M1_U4_U1_or2_inv_1__20_)
         );
  INVXL U25033 ( .A(M1_U4_U1_enc_tree_1__1__12_), .Y(M1_U4_U1_or2_inv_1__12_)
         );
  INVXL U25034 ( .A(M1_U3_U1_enc_tree_1__1__28_), .Y(M1_U3_U1_or2_inv_1__28_)
         );
  INVXL U25035 ( .A(M1_U3_U1_or2_tree_1__2__24_), .Y(M1_U3_U1_or2_inv_1__24_)
         );
  INVXL U25036 ( .A(M1_U3_U1_enc_tree_1__1__20_), .Y(M1_U3_U1_or2_inv_1__20_)
         );
  INVXL U25037 ( .A(M1_U3_U1_enc_tree_1__1__12_), .Y(M1_U3_U1_or2_inv_1__12_)
         );
  NAND4XL U25038 ( .A(n23181), .B(n23180), .C(n23179), .D(n23178), .Y(n23187)
         );
  NAND4XL U25039 ( .A(n23185), .B(n23184), .C(n23183), .D(n23182), .Y(n23186)
         );
  NOR2XL U25040 ( .A(n23187), .B(n23186), .Y(n23188) );
  AOI2BB1XL U25041 ( .A0N(n23189), .A1N(n23188), .B0(n9027), .Y(n23190) );
  NOR3X1 U25042 ( .A(n23192), .B(n23191), .C(n23190), .Y(n25697) );
  AOI21XL U25043 ( .A0(n5604), .A1(n26048), .B0(n23194), .Y(n23195) );
  NAND4XL U25044 ( .A(n23206), .B(n23205), .C(n23204), .D(n23203), .Y(n23212)
         );
  NAND4XL U25045 ( .A(n23210), .B(n23209), .C(n23208), .D(n23207), .Y(n23211)
         );
  NOR2XL U25046 ( .A(n23212), .B(n23211), .Y(n23213) );
  CMPR22X1 U25047 ( .A(n23218), .B(n23217), .CO(M6_mult_x_15_n727), .S(n10885)
         );
  INVXL U25048 ( .A(M5_U3_U1_enc_tree_1__1__20_), .Y(M5_U3_U1_or2_inv_1__20_)
         );
  INVXL U25049 ( .A(M5_U3_U1_enc_tree_1__1__12_), .Y(M5_U3_U1_or2_inv_1__12_)
         );
  INVXL U25050 ( .A(M5_U3_U1_or2_tree_0__1__28_), .Y(M5_U3_U1_or2_inv_0__28_)
         );
  INVXL U25051 ( .A(M5_U3_U1_or2_tree_0__1__20_), .Y(M5_U3_U1_or2_inv_0__20_)
         );
  INVXL U25052 ( .A(M0_U3_U1_enc_tree_1__1__28_), .Y(M0_U3_U1_or2_inv_1__28_)
         );
  INVXL U25053 ( .A(M0_U3_U1_enc_tree_1__1__20_), .Y(M0_U3_U1_or2_inv_1__20_)
         );
  INVXL U25054 ( .A(M0_U3_U1_enc_tree_1__1__12_), .Y(M0_U3_U1_or2_inv_1__12_)
         );
  INVXL U25055 ( .A(M0_U4_U1_enc_tree_1__1__20_), .Y(M0_U4_U1_or2_inv_1__20_)
         );
  INVXL U25056 ( .A(M0_U4_U1_enc_tree_1__1__12_), .Y(M0_U4_U1_or2_inv_1__12_)
         );
  INVXL U25057 ( .A(M0_U3_U1_or2_tree_0__1__28_), .Y(M0_U3_U1_or2_inv_0__28_)
         );
  INVXL U25058 ( .A(M0_U3_U1_or2_tree_0__1__20_), .Y(M0_U3_U1_or2_inv_0__20_)
         );
  INVXL U25059 ( .A(M0_b_5_), .Y(M0_U4_U1_or2_inv_0__26_) );
  INVXL U25060 ( .A(M0_b_9_), .Y(M0_U4_U1_or2_inv_0__22_) );
  INVXL U25061 ( .A(M0_U4_U1_or2_tree_0__1__20_), .Y(M0_U4_U1_or2_inv_0__20_)
         );
  INVXL U25062 ( .A(M0_b_13_), .Y(M0_U4_U1_or2_inv_0__18_) );
  INVXL U25063 ( .A(M0_b_17_), .Y(M0_U4_U1_or2_inv_0__14_) );
  INVXL U25064 ( .A(M0_b_21_), .Y(M0_U4_U1_or2_inv_0__10_) );
  INVXL U25065 ( .A(M3_U3_U1_enc_tree_1__1__20_), .Y(M3_U3_U1_or2_inv_1__20_)
         );
  INVXL U25066 ( .A(M3_U3_U1_enc_tree_1__1__12_), .Y(M3_U3_U1_or2_inv_1__12_)
         );
  INVXL U25067 ( .A(M3_U3_U1_or2_tree_0__1__28_), .Y(M3_U3_U1_or2_inv_0__28_)
         );
  INVXL U25068 ( .A(M3_U3_U1_or2_tree_0__1__20_), .Y(M3_U3_U1_or2_inv_0__20_)
         );
  INVXL U25069 ( .A(M4_U3_U1_enc_tree_1__1__28_), .Y(M4_U3_U1_or2_inv_1__28_)
         );
  INVXL U25070 ( .A(M4_U3_U1_or2_tree_1__2__24_), .Y(M4_U3_U1_or2_inv_1__24_)
         );
  INVXL U25071 ( .A(M4_U3_U1_enc_tree_1__1__20_), .Y(M4_U3_U1_or2_inv_1__20_)
         );
  INVXL U25072 ( .A(M4_U3_U1_enc_tree_1__1__12_), .Y(M4_U3_U1_or2_inv_1__12_)
         );
  INVXL U25073 ( .A(M4_U3_U1_or2_tree_0__1__28_), .Y(M4_U3_U1_or2_inv_0__28_)
         );
  INVXL U25074 ( .A(M4_U3_U1_or2_tree_0__2__24_), .Y(M4_U3_U1_or2_inv_0__24_)
         );
  INVXL U25075 ( .A(M4_U3_U1_or2_tree_0__1__20_), .Y(M4_U3_U1_or2_inv_0__20_)
         );
  INVXL U25076 ( .A(M4_U4_U1_or2_tree_0__1__20_), .Y(M3_U4_U1_or2_inv_0__20_)
         );
  INVXL U25077 ( .A(M2_U4_U1_or2_tree_0__1__28_), .Y(M2_U4_U1_or2_inv_0__28_)
         );
  INVXL U25078 ( .A(M2_U4_U1_or2_tree_0__2__24_), .Y(M2_U4_U1_or2_inv_0__24_)
         );
  INVXL U25079 ( .A(M2_U4_U1_or2_tree_0__1__20_), .Y(M2_U4_U1_or2_inv_0__20_)
         );
  INVXL U25080 ( .A(M2_b_13_), .Y(M2_U4_U1_or2_inv_0__18_) );
  INVXL U25081 ( .A(n23222), .Y(M2_U4_U1_or2_inv_0__10_) );
  INVXL U25082 ( .A(M2_U3_U1_or2_tree_0__1__28_), .Y(M2_U3_U1_or2_inv_0__28_)
         );
  INVXL U25083 ( .A(M2_U3_U1_or2_tree_0__2__24_), .Y(M2_U3_U1_or2_inv_0__24_)
         );
  INVXL U25084 ( .A(M2_U3_U1_or2_tree_0__1__20_), .Y(M2_U3_U1_or2_inv_0__20_)
         );
  INVXL U25085 ( .A(M2_U4_U1_enc_tree_1__1__28_), .Y(M2_U4_U1_or2_inv_1__28_)
         );
  INVXL U25086 ( .A(M2_U4_U1_or2_tree_1__2__24_), .Y(M2_U4_U1_or2_inv_1__24_)
         );
  INVXL U25087 ( .A(M2_U4_U1_enc_tree_1__1__20_), .Y(M2_U4_U1_or2_inv_1__20_)
         );
  INVXL U25088 ( .A(M2_U4_U1_enc_tree_1__1__12_), .Y(M2_U4_U1_or2_inv_1__12_)
         );
  INVXL U25089 ( .A(M2_U3_U1_enc_tree_1__1__28_), .Y(M2_U3_U1_or2_inv_1__28_)
         );
  INVXL U25090 ( .A(M2_U3_U1_or2_tree_1__2__24_), .Y(M2_U3_U1_or2_inv_1__24_)
         );
  INVXL U25091 ( .A(M2_U3_U1_enc_tree_1__1__20_), .Y(M2_U3_U1_or2_inv_1__20_)
         );
  INVXL U25092 ( .A(M2_U3_U1_enc_tree_1__2__12_), .Y(
        M2_U3_U1_enc_tree_1__3__8_) );
  INVXL U25093 ( .A(M2_U3_U1_enc_tree_1__1__12_), .Y(M2_U3_U1_or2_inv_1__12_)
         );
  INVXL U25094 ( .A(M2_U3_U1_enc_tree_2__2__24_), .Y(M2_U3_U1_or2_inv_2__24_)
         );
  INVXL U25095 ( .A(M2_U4_U1_enc_tree_2__2__24_), .Y(M2_U4_U1_or2_inv_2__24_)
         );
  NOR2X2 U25096 ( .A(n4767), .B(n23228), .Y(n23419) );
  AOI222XL U25097 ( .A0(n23234), .A1(n3216), .B0(n3023), .B1(w1[283]), .C0(
        n3061), .C1(w1[315]), .Y(n2119) );
  AOI222XL U25098 ( .A0(n23248), .A1(n25541), .B0(w1[265]), .B1(n4577), .C0(
        n3061), .C1(w1[297]), .Y(n2047) );
  AOI222XL U25099 ( .A0(n23249), .A1(n3216), .B0(w1[266]), .B1(n4577), .C0(
        n23088), .C1(w1[298]), .Y(n2051) );
  AOI21XL U25100 ( .A0(n23324), .A1(n23429), .B0(n23253), .Y(n23254) );
  XNOR2XL U25101 ( .A(n23273), .B(n23272), .Y(n23274) );
  NAND2XL U25102 ( .A(n23346), .B(n23318), .Y(n23320) );
  AOI222XL U25103 ( .A0(n23325), .A1(n3216), .B0(w1[260]), .B1(n4578), .C0(
        n3061), .C1(w1[292]), .Y(n2027) );
  NOR2XL U25104 ( .A(n23330), .B(n23329), .Y(n23331) );
  AOI222XL U25105 ( .A0(n23352), .A1(n3216), .B0(w1[264]), .B1(n4577), .C0(
        n23088), .C1(w1[296]), .Y(n2043) );
  AOI222XL U25106 ( .A0(n23353), .A1(n21112), .B0(w1[262]), .B1(n4576), .C0(
        n23088), .C1(w1[294]), .Y(n2035) );
  AOI222XL U25107 ( .A0(n23354), .A1(n3216), .B0(w1[261]), .B1(n4578), .C0(
        n3061), .C1(w1[293]), .Y(n2031) );
  AOI222XL U25108 ( .A0(n23356), .A1(n3216), .B0(w1[256]), .B1(n4578), .C0(
        n23088), .C1(w1[288]), .Y(n2011) );
  AOI222XL U25109 ( .A0(n23357), .A1(n21112), .B0(w1[263]), .B1(n4577), .C0(
        n3061), .C1(w1[295]), .Y(n2039) );
  AOI222XL U25110 ( .A0(n23358), .A1(n3216), .B0(w1[273]), .B1(n4576), .C0(
        n23088), .C1(w1[305]), .Y(n2079) );
  AOI222XL U25111 ( .A0(n23359), .A1(n3216), .B0(w1[271]), .B1(n4577), .C0(
        n3061), .C1(w1[303]), .Y(n2071) );
  AOI222XL U25112 ( .A0(n23360), .A1(n25541), .B0(w1[268]), .B1(n4577), .C0(
        n23088), .C1(w1[300]), .Y(n2059) );
  AOI222XL U25113 ( .A0(n23361), .A1(n25541), .B0(w1[267]), .B1(n4577), .C0(
        n23088), .C1(w1[299]), .Y(n2055) );
  AOI222XL U25114 ( .A0(n23362), .A1(n3216), .B0(w1[274]), .B1(n4577), .C0(
        n23088), .C1(w1[306]), .Y(n2083) );
  AOI222XL U25115 ( .A0(n23363), .A1(n25541), .B0(w1[257]), .B1(n4578), .C0(
        n3061), .C1(w1[289]), .Y(n2015) );
  AOI222XL U25116 ( .A0(n23364), .A1(n25541), .B0(w1[258]), .B1(n4578), .C0(
        n3061), .C1(w1[290]), .Y(n2019) );
  AOI222XL U25117 ( .A0(n23365), .A1(n25541), .B0(w1[259]), .B1(n4577), .C0(
        n23088), .C1(w1[291]), .Y(n2023) );
  AOI222XL U25118 ( .A0(n23366), .A1(n3216), .B0(w1[272]), .B1(n4577), .C0(
        n3061), .C1(w1[304]), .Y(n2075) );
  AOI222XL U25119 ( .A0(n23367), .A1(n25541), .B0(w1[270]), .B1(n4576), .C0(
        n3061), .C1(w1[302]), .Y(n2067) );
  AOI222XL U25120 ( .A0(n23368), .A1(n25541), .B0(w1[269]), .B1(n4577), .C0(
        n23088), .C1(w1[301]), .Y(n2063) );
  NAND2XL U25121 ( .A(n23383), .B(n23376), .Y(n23378) );
  AOI222XL U25122 ( .A0(n23389), .A1(n3216), .B0(w1[276]), .B1(n4576), .C0(
        n3061), .C1(w1[308]), .Y(n2091) );
  AOI222XL U25123 ( .A0(n23390), .A1(n3216), .B0(w1[275]), .B1(n4576), .C0(
        n23088), .C1(w1[307]), .Y(n2087) );
  AOI222XL U25124 ( .A0(n23391), .A1(n3216), .B0(w1[277]), .B1(n4576), .C0(
        n23088), .C1(w1[309]), .Y(n2095) );
  AOI222X1 U25125 ( .A0(n23394), .A1(n23419), .B0(n23418), .B1(n23393), .C0(
        n23392), .C1(n23415), .Y(n23395) );
  INVX1 U25126 ( .A(n23395), .Y(n23424) );
  AOI222X1 U25127 ( .A0(n23398), .A1(n23419), .B0(n23418), .B1(n23397), .C0(
        n23396), .C1(n23415), .Y(n23399) );
  INVX1 U25128 ( .A(n23399), .Y(n23423) );
  AOI222X1 U25129 ( .A0(n23402), .A1(n23419), .B0(n23418), .B1(n23401), .C0(
        n23400), .C1(n23415), .Y(n23403) );
  INVX1 U25130 ( .A(n23403), .Y(n23430) );
  AOI222X1 U25131 ( .A0(n23406), .A1(n23419), .B0(n23418), .B1(n23405), .C0(
        n23404), .C1(n23415), .Y(n23407) );
  INVX1 U25132 ( .A(n23407), .Y(n23422) );
  AOI222X1 U25133 ( .A0(n23409), .A1(n23419), .B0(n23418), .B1(n22222), .C0(
        n23408), .C1(n23415), .Y(n23410) );
  INVX1 U25134 ( .A(n23410), .Y(n23425) );
  INVX1 U25135 ( .A(n23414), .Y(n23426) );
  AOI222X1 U25136 ( .A0(n23420), .A1(n23419), .B0(n23418), .B1(n23417), .C0(
        n23416), .C1(n23415), .Y(n23421) );
  INVX1 U25137 ( .A(n23421), .Y(n23427) );
  NOR2XL U25138 ( .A(n23431), .B(n23442), .Y(n23432) );
  NAND2XL U25139 ( .A(n23744), .B(n23432), .Y(n23434) );
  XOR2X1 U25140 ( .A(n23434), .B(n23433), .Y(n23631) );
  INVXL U25141 ( .A(n23436), .Y(n23438) );
  NAND2XL U25142 ( .A(n23438), .B(n23437), .Y(n23439) );
  XOR2X1 U25143 ( .A(n23486), .B(n23439), .Y(n25294) );
  NAND2XL U25144 ( .A(n25298), .B(n23794), .Y(n23440) );
  NAND2XL U25145 ( .A(n23744), .B(n3141), .Y(n23443) );
  XOR2X1 U25146 ( .A(n23443), .B(n23442), .Y(n23630) );
  NAND2XL U25147 ( .A(n23744), .B(n23446), .Y(n23449) );
  INVXL U25148 ( .A(n23447), .Y(n23448) );
  XOR2X1 U25149 ( .A(n23449), .B(n23448), .Y(n23880) );
  AOI22X1 U25150 ( .A0(n3081), .A1(n23630), .B0(n23880), .B1(n4267), .Y(n24155) );
  XOR2X1 U25151 ( .A(n23451), .B(n5410), .Y(n24169) );
  AOI22XL U25152 ( .A0(n24169), .A1(n23794), .B0(n2983), .B1(temp1[9]), .Y(
        n23453) );
  NAND2XL U25153 ( .A(n24160), .B(n23795), .Y(n23452) );
  OAI211XL U25154 ( .A0(n24155), .A1(n4583), .B0(n23453), .C0(n23452), .Y(
        n2545) );
  INVX1 U25155 ( .A(n23458), .Y(n23459) );
  NAND2X1 U25156 ( .A(n23734), .B(n23527), .Y(n23461) );
  XOR2X1 U25157 ( .A(n23461), .B(n3033), .Y(n25553) );
  AOI22XL U25158 ( .A0(n23949), .A1(n23885), .B0(n23947), .B1(n23726), .Y(
        n23471) );
  INVXL U25159 ( .A(n23476), .Y(n23477) );
  AOI22X1 U25160 ( .A0(n23483), .A1(n23883), .B0(n5211), .B1(n6199), .Y(n24460) );
  AOI22XL U25161 ( .A0(n23794), .A1(n25294), .B0(n2984), .B1(temp1[0]), .Y(
        n23488) );
  NAND2XL U25162 ( .A(n23795), .B(n25335), .Y(n23487) );
  OAI211XL U25163 ( .A0(n24460), .A1(n4583), .B0(n23488), .C0(n23487), .Y(
        n2554) );
  NAND2X1 U25164 ( .A(n3132), .B(n23489), .Y(n23490) );
  INVXL U25165 ( .A(n23491), .Y(n23493) );
  NAND2XL U25166 ( .A(n23493), .B(n23492), .Y(n23531) );
  XOR2X1 U25167 ( .A(n23511), .B(n23733), .Y(n25503) );
  NAND2XL U25168 ( .A(n23527), .B(n23512), .Y(n23523) );
  INVXL U25169 ( .A(n23513), .Y(n23525) );
  NOR2XL U25170 ( .A(n23523), .B(n23525), .Y(n23514) );
  XOR2X1 U25171 ( .A(n23517), .B(n23516), .Y(n25527) );
  NAND2XL U25172 ( .A(n23734), .B(n23518), .Y(n23520) );
  INVXL U25173 ( .A(n23523), .Y(n23524) );
  NAND2XL U25174 ( .A(n23734), .B(n23524), .Y(n23526) );
  XOR2X1 U25175 ( .A(n23526), .B(n23525), .Y(n25528) );
  INVXL U25176 ( .A(n23531), .Y(n23532) );
  AOI22XL U25177 ( .A0(n23939), .A1(n23949), .B0(n23544), .B1(n23947), .Y(
        n23545) );
  INVXL U25178 ( .A(n23551), .Y(n23552) );
  XOR2X1 U25179 ( .A(n23553), .B(n23552), .Y(n25762) );
  NAND2XL U25180 ( .A(n25762), .B(n25636), .Y(n23554) );
  OAI211XL U25181 ( .A0(n25747), .A1(n4586), .B0(n23555), .C0(n23554), .Y(
        n2573) );
  NOR2X1 U25182 ( .A(n5033), .B(n5465), .Y(n23557) );
  AOI22XL U25183 ( .A0(n24206), .A1(n25638), .B0(n2983), .B1(temp2[16]), .Y(
        n23560) );
  NAND2XL U25184 ( .A(n25636), .B(n24218), .Y(n23559) );
  OAI211XL U25185 ( .A0(n24821), .A1(n4583), .B0(n23560), .C0(n23559), .Y(
        n2585) );
  NAND2XL U25186 ( .A(n4643), .B(n23561), .Y(n23562) );
  XOR2X1 U25187 ( .A(n23562), .B(n24253), .Y(n25635) );
  AOI22XL U25188 ( .A0(n25638), .A1(n25635), .B0(n2984), .B1(temp2[1]), .Y(
        n23564) );
  NAND2XL U25189 ( .A(n24057), .B(n25636), .Y(n23563) );
  NAND2XL U25190 ( .A(n24244), .B(n25638), .Y(n23566) );
  OAI211XL U25191 ( .A0(n24913), .A1(n4586), .B0(n23567), .C0(n23566), .Y(
        n2579) );
  AOI22XL U25192 ( .A0(n24140), .A1(n23794), .B0(n2983), .B1(temp1[5]), .Y(
        n23571) );
  NAND2XL U25193 ( .A(n24135), .B(n23795), .Y(n23570) );
  AOI22XL U25194 ( .A0(n24192), .A1(n23794), .B0(n2984), .B1(temp1[12]), .Y(
        n23575) );
  NAND2XL U25195 ( .A(n24183), .B(n23795), .Y(n23574) );
  OAI211XL U25196 ( .A0(n24177), .A1(n4584), .B0(n23575), .C0(n23574), .Y(
        n2542) );
  CLKINVX3 U25197 ( .A(n23764), .Y(n24739) );
  CLKINVX3 U25198 ( .A(n20748), .Y(n25656) );
  OAI21XL U25199 ( .A0(n23577), .A1(n3057), .B0(n23576), .Y(n23578) );
  INVXL U25200 ( .A(n23583), .Y(n23581) );
  CLKINVX3 U25201 ( .A(n23764), .Y(n25815) );
  OAI21XL U25202 ( .A0(n23768), .A1(n3057), .B0(n23584), .Y(n23585) );
  AOI21XL U25203 ( .A0(n23769), .A1(n25675), .B0(n23585), .Y(n2408) );
  AOI22XL U25204 ( .A0(n24206), .A1(n25636), .B0(n2984), .B1(temp2[15]), .Y(
        n23587) );
  NAND2XL U25205 ( .A(n24210), .B(n25638), .Y(n23586) );
  OAI211XL U25206 ( .A0(n24769), .A1(n4584), .B0(n23587), .C0(n23586), .Y(
        n2587) );
  AOI22XL U25207 ( .A0(n23949), .A1(n23899), .B0(n23947), .B1(n23907), .Y(
        n23602) );
  NAND2XL U25208 ( .A(n23829), .B(n23754), .Y(n23606) );
  XOR2X1 U25209 ( .A(n23606), .B(n23605), .Y(n23607) );
  CLKINVX3 U25210 ( .A(n23764), .Y(n25025) );
  OAI21XL U25211 ( .A0(n23720), .A1(n3057), .B0(n23609), .Y(n23610) );
  AOI21XL U25212 ( .A0(n23721), .A1(n3060), .B0(n23610), .Y(n2426) );
  INVXL U25213 ( .A(n23827), .Y(n23613) );
  NAND2XL U25214 ( .A(n23829), .B(n23613), .Y(n23614) );
  XOR2X1 U25215 ( .A(n23614), .B(n23826), .Y(n23615) );
  OAI21XL U25216 ( .A0(n25323), .A1(n3057), .B0(n23617), .Y(n23618) );
  AOI21XL U25217 ( .A0(n25733), .A1(n6161), .B0(n23618), .Y(n2428) );
  NOR2XL U25218 ( .A(n24562), .B(n23621), .Y(n23623) );
  INVXL U25219 ( .A(n23625), .Y(n23622) );
  AOI222XL U25220 ( .A0(n24548), .A1(n25744), .B0(n25743), .B1(y20[5]), .C0(
        n25568), .C1(n20890), .Y(n2365) );
  AOI22XL U25221 ( .A0(n24127), .A1(n23794), .B0(n2983), .B1(temp1[3]), .Y(
        n23629) );
  NAND2XL U25222 ( .A(n24123), .B(n23795), .Y(n23628) );
  OAI211XL U25223 ( .A0(n24491), .A1(n4581), .B0(n23629), .C0(n23628), .Y(
        n2551) );
  NAND2XL U25224 ( .A(n24174), .B(n23794), .Y(n23632) );
  INVX1 U25225 ( .A(n23639), .Y(n23633) );
  OAI2BB1X1 U25226 ( .A0N(n24360), .A1N(n23643), .B0(n23647), .Y(mul5_out[24])
         );
  NAND2XL U25227 ( .A(n23744), .B(n3083), .Y(n23649) );
  NAND2XL U25228 ( .A(n3895), .B(n3894), .Y(n23652) );
  XOR2X1 U25229 ( .A(n23651), .B(n23652), .Y(n24201) );
  AOI22XL U25230 ( .A0(n24201), .A1(n23794), .B0(n2983), .B1(temp1[13]), .Y(
        n23654) );
  NAND2XL U25231 ( .A(n24192), .B(n23795), .Y(n23653) );
  OAI21XL U25232 ( .A0(n23656), .A1(n3057), .B0(n23655), .Y(n23657) );
  AOI21XL U25233 ( .A0(n23658), .A1(n6161), .B0(n23657), .Y(n2414) );
  ADDHXL U25234 ( .A(n23660), .B(n23661), .CO(n23663), .S(n20801) );
  INVXL U25235 ( .A(n23669), .Y(n23671) );
  INVXL U25236 ( .A(n25245), .Y(n23670) );
  OAI21XL U25237 ( .A0(n23674), .A1(n23671), .B0(n23670), .Y(n23672) );
  OAI21XL U25238 ( .A0(n23678), .A1(n23677), .B0(n23715), .Y(n23679) );
  AOI22XL U25239 ( .A0(n23681), .A1(n3223), .B0(n25723), .B1(temp0[30]), .Y(
        n23688) );
  NAND2XL U25240 ( .A(n23839), .B(n3065), .Y(n23687) );
  OAI211XL U25241 ( .A0(n25851), .A1(n3121), .B0(n23688), .C0(n23687), .Y(
        n2556) );
  AOI22XL U25242 ( .A0(n23873), .A1(n23691), .B0(n23871), .B1(n23690), .Y(
        n23692) );
  INVXL U25243 ( .A(n25801), .Y(n23695) );
  AOI21XL U25244 ( .A0(n23839), .A1(n3060), .B0(n23696), .Y(n2452) );
  INVXL U25245 ( .A(n23697), .Y(mul5_out[6]) );
  OAI21XL U25246 ( .A0(n23699), .A1(n3057), .B0(n23698), .Y(n23700) );
  AOI21XL U25247 ( .A0(n23701), .A1(n24525), .B0(n23700), .Y(n2406) );
  AOI22XL U25248 ( .A0(n24227), .A1(n23794), .B0(n2984), .B1(temp1[16]), .Y(
        n23705) );
  NAND2XL U25249 ( .A(n24220), .B(n23795), .Y(n23704) );
  OAI211XL U25250 ( .A0(n24847), .A1(n4586), .B0(n23714), .C0(n23713), .Y(
        n2536) );
  INVXL U25251 ( .A(n23862), .Y(n23718) );
  AOI22XL U25252 ( .A0(n23949), .A1(n23726), .B0(n23947), .B1(n23725), .Y(
        n23727) );
  NAND2XL U25253 ( .A(n23737), .B(n23738), .Y(n23740) );
  INVXL U25254 ( .A(n23745), .Y(n23746) );
  INVXL U25255 ( .A(n23749), .Y(n23750) );
  OAI21XL U25256 ( .A0(n23756), .A1(n3057), .B0(n23755), .Y(n23757) );
  AOI21XL U25257 ( .A0(n23758), .A1(n25675), .B0(n23757), .Y(n2424) );
  AOI22XL U25258 ( .A0(n23873), .A1(n23761), .B0(n23871), .B1(n23760), .Y(
        n23762) );
  OAI21X1 U25259 ( .A0(n4788), .A1(n23763), .B0(n23762), .Y(n24321) );
  INVXL U25260 ( .A(n24321), .Y(n23766) );
  AOI22XL U25261 ( .A0(n24739), .A1(y10[23]), .B0(n3122), .B1(y12[23]), .Y(
        n23765) );
  AOI21XL U25262 ( .A0(n23972), .A1(n3060), .B0(n23767), .Y(n2438) );
  INVXL U25263 ( .A(n23773), .Y(n23771) );
  XNOR2XL U25264 ( .A(n23771), .B(n25301), .Y(n23772) );
  AOI22X1 U25265 ( .A0(n20385), .A1(n23773), .B0(n25300), .B1(n23772), .Y(
        n24473) );
  AOI222XL U25266 ( .A0(n24475), .A1(n25744), .B0(n25743), .B1(y20[1]), .C0(
        n25624), .C1(n20890), .Y(n2361) );
  INVXL U25267 ( .A(n23777), .Y(n23778) );
  OAI21XL U25268 ( .A0(n25703), .A1(n25700), .B0(n23786), .Y(n23788) );
  OR3XL U25269 ( .A(n25832), .B(n23786), .C(n23785), .Y(n23787) );
  AOI22XL U25270 ( .A0(n23794), .A1(n24211), .B0(n2984), .B1(temp1[14]), .Y(
        n23797) );
  NAND2XL U25271 ( .A(n24201), .B(n23795), .Y(n23796) );
  OAI211XL U25272 ( .A0(n24715), .A1(n4583), .B0(n23797), .C0(n23796), .Y(
        n2540) );
  INVXL U25273 ( .A(n23798), .Y(n23800) );
  NOR2XL U25274 ( .A(n23800), .B(n23799), .Y(n23801) );
  NAND2XL U25275 ( .A(n23829), .B(n23801), .Y(n23803) );
  AOI22XL U25276 ( .A0(n23873), .A1(n23811), .B0(n23871), .B1(n23810), .Y(
        n23812) );
  CLKINVX3 U25277 ( .A(n25292), .Y(n25711) );
  AOI222XL U25278 ( .A0(n24421), .A1(n3216), .B0(w1[313]), .B1(n4576), .C0(
        n3061), .C1(w1[345]), .Y(n2108) );
  AOI22XL U25279 ( .A0(n23873), .A1(n23817), .B0(n23871), .B1(n23816), .Y(
        n23818) );
  AOI222XL U25280 ( .A0(n25720), .A1(n25744), .B0(y20[26]), .B1(n25743), .C0(
        n24417), .C1(n20890), .Y(n2386) );
  NOR2XL U25281 ( .A(n23827), .B(n23826), .Y(n23828) );
  NAND2XL U25282 ( .A(n23829), .B(n23828), .Y(n23831) );
  OAI21XL U25283 ( .A0(n23836), .A1(n3057), .B0(n23834), .Y(n23835) );
  AOI21XL U25284 ( .A0(n23837), .A1(n6161), .B0(n23835), .Y(n2430) );
  AOI222XL U25285 ( .A0(n23839), .A1(n25737), .B0(y20[30]), .B1(n25743), .C0(
        n25801), .C1(n20890), .Y(n2390) );
  OAI21XL U25286 ( .A0(n23841), .A1(n3057), .B0(n23840), .Y(n23842) );
  INVXL U25287 ( .A(n23843), .Y(n23847) );
  AOI22XL U25288 ( .A0(n23873), .A1(n23845), .B0(n23871), .B1(n23844), .Y(
        n23846) );
  OAI21X1 U25289 ( .A0(n4788), .A1(n23847), .B0(n23846), .Y(n25683) );
  ADDHXL U25290 ( .A(n23850), .B(n23849), .CO(n23684), .S(n23852) );
  AOI21XL U25291 ( .A0(n23850), .A1(n23864), .B0(n23863), .Y(n23851) );
  AOI222XL U25292 ( .A0(n25840), .A1(n25737), .B0(y20[29]), .B1(n25743), .C0(
        n25683), .C1(n20890), .Y(n2389) );
  AOI222XL U25293 ( .A0(n24447), .A1(n25744), .B0(y20[28]), .B1(n25743), .C0(
        n24451), .C1(n20890), .Y(n2388) );
  AOI222XL U25294 ( .A0(n24451), .A1(n3216), .B0(w1[316]), .B1(n4578), .C0(
        n23088), .C1(w1[348]), .Y(n2120) );
  AOI21XL U25295 ( .A0(n23854), .A1(n23864), .B0(n23863), .Y(n23855) );
  AOI22XL U25296 ( .A0(n23873), .A1(n23859), .B0(n23871), .B1(n23858), .Y(
        n23860) );
  OAI21X1 U25297 ( .A0(n4788), .A1(n23861), .B0(n23860), .Y(n25080) );
  AOI222XL U25298 ( .A0(n25076), .A1(n25737), .B0(y20[27]), .B1(n25743), .C0(
        n25080), .C1(n20890), .Y(n2387) );
  ADDHXL U25299 ( .A(n23865), .B(n23862), .CO(n23781), .S(n23867) );
  AOI21XL U25300 ( .A0(n23865), .A1(n23864), .B0(n23863), .Y(n23866) );
  AOI22XL U25301 ( .A0(n23873), .A1(n23872), .B0(n23871), .B1(n23870), .Y(
        n23874) );
  INVXL U25302 ( .A(n25712), .Y(n23877) );
  AOI21XL U25303 ( .A0(n25707), .A1(n24525), .B0(n23878), .Y(n2440) );
  AOI222XL U25304 ( .A0(n25707), .A1(n25744), .B0(y20[24]), .B1(n25743), .C0(
        n25712), .C1(n20890), .Y(n2384) );
  AOI22X1 U25305 ( .A0(n3081), .A1(n23880), .B0(n23879), .B1(n5211), .Y(n24595) );
  AOI22X2 U25306 ( .A0(n3081), .A1(n23882), .B0(n23881), .B1(n4267), .Y(n24888) );
  AOI22XL U25307 ( .A0(n23949), .A1(n23886), .B0(n23947), .B1(n23885), .Y(
        n23887) );
  AOI22XL U25308 ( .A0(n23932), .A1(n23949), .B0(n23947), .B1(n23899), .Y(
        n23900) );
  AOI22XL U25309 ( .A0(n23949), .A1(n23907), .B0(n23947), .B1(n23948), .Y(
        n23908) );
  AOI22XL U25310 ( .A0(n23949), .A1(n23927), .B0(n23947), .B1(n23919), .Y(
        n23920) );
  AOI22XL U25311 ( .A0(n23949), .A1(n23928), .B0(n23947), .B1(n23927), .Y(
        n23929) );
  AOI22XL U25312 ( .A0(n23933), .A1(n23949), .B0(n23947), .B1(n23932), .Y(
        n23934) );
  AOI22XL U25313 ( .A0(n23940), .A1(n23949), .B0(n23947), .B1(n23939), .Y(
        n23941) );
  INVXL U25314 ( .A(n23961), .Y(n23958) );
  AOI222X1 U25315 ( .A0(n23966), .A1(n24430), .B0(n24427), .B1(n23965), .C0(
        n23964), .C1(n24428), .Y(n24317) );
  AOI222XL U25316 ( .A0(n24325), .A1(n4710), .B0(in_valid_w2), .B1(weight2[23]), .C0(w2[87]), .C1(n25822), .Y(n2223) );
  OAI21XL U25317 ( .A0(n3061), .A1(n23967), .B0(n3024), .Y(n23968) );
  AOI21XL U25318 ( .A0(n23970), .A1(n23969), .B0(n23968), .Y(n2490) );
  AOI222XL U25319 ( .A0(n23972), .A1(n25744), .B0(y20[23]), .B1(n25743), .C0(
        n24321), .C1(n20890), .Y(n2383) );
  MXI2XL U25320 ( .A(n23974), .B(n23973), .S0(n3057), .Y(N42) );
  NAND2XL U25321 ( .A(n3057), .B(valid[2]), .Y(n23975) );
  OAI21XL U25322 ( .A0(n23973), .A1(n3057), .B0(n23975), .Y(N41) );
  NAND2XL U25323 ( .A(n24011), .B(n23976), .Y(n24013) );
  AOI21XL U25324 ( .A0(n23978), .A1(n23977), .B0(n24012), .Y(n23979) );
  INVXL U25325 ( .A(n23979), .Y(n24009) );
  NOR3XL U25326 ( .A(learning_rate[25]), .B(learning_rate[26]), .C(
        learning_rate[28]), .Y(n23981) );
  NAND4XL U25327 ( .A(learning_rate[23]), .B(n23982), .C(n23981), .D(n23980), 
        .Y(n23983) );
  NOR3BXL U25328 ( .AN(n24013), .B(n24009), .C(n23983), .Y(n23984) );
  OAI21XL U25329 ( .A0(n23987), .A1(n23988), .B0(n23997), .Y(n2633) );
  OAI21XL U25330 ( .A0(n23987), .A1(n23989), .B0(n23997), .Y(n2634) );
  OAI21XL U25331 ( .A0(n23987), .A1(n23990), .B0(n23997), .Y(n2638) );
  OAI21XL U25332 ( .A0(n23987), .A1(n23991), .B0(n23997), .Y(n2639) );
  OAI21XL U25333 ( .A0(n23987), .A1(n23992), .B0(n23997), .Y(n2641) );
  OAI21XL U25334 ( .A0(n23987), .A1(n23993), .B0(n23997), .Y(n2642) );
  OAI21XL U25335 ( .A0(n23987), .A1(n23994), .B0(n23997), .Y(n2643) );
  OAI21XL U25336 ( .A0(n23987), .A1(n23995), .B0(n23997), .Y(n2644) );
  OAI21XL U25337 ( .A0(n23987), .A1(n23996), .B0(n23997), .Y(n2646) );
  OAI21XL U25338 ( .A0(n23987), .A1(n23998), .B0(n23997), .Y(n2647) );
  OAI21XL U25339 ( .A0(n23987), .A1(n23999), .B0(n23997), .Y(n2648) );
  OAI21XL U25340 ( .A0(n23987), .A1(n24000), .B0(n23997), .Y(n2649) );
  OAI21XL U25341 ( .A0(n23987), .A1(n24001), .B0(n23997), .Y(n2651) );
  OAI21XL U25342 ( .A0(n24003), .A1(n24006), .B0(n24002), .Y(n24004) );
  OAI21XL U25343 ( .A0(n25856), .A1(n24006), .B0(n24005), .Y(n2626) );
  INVXL U25344 ( .A(learning_rate[30]), .Y(n24017) );
  OAI21XL U25345 ( .A0(n24013), .A1(n24012), .B0(n24011), .Y(n24014) );
  NAND2XL U25346 ( .A(n24015), .B(n24014), .Y(n24016) );
  OAI21XL U25347 ( .A0(n25856), .A1(n24017), .B0(n24016), .Y(n2621) );
  AOI222XL U25348 ( .A0(n25845), .A1(n25292), .B0(weight2[30]), .B1(
        in_valid_w2), .C0(w2[94]), .C1(n25822), .Y(n2230) );
  AOI21XL U25349 ( .A0(data[126]), .A1(n4584), .B0(n24021), .Y(n1740) );
  AOI21XL U25350 ( .A0(data[119]), .A1(n4585), .B0(n24023), .Y(n1733) );
  AOI21XL U25351 ( .A0(data[118]), .A1(n4583), .B0(n24024), .Y(n1732) );
  NAND2XL U25352 ( .A(n24031), .B(n25774), .Y(n24039) );
  INVX2 U25353 ( .A(n24035), .Y(n24031) );
  NAND2XL U25354 ( .A(n25778), .B(n24032), .Y(n24038) );
  OAI21X2 U25355 ( .A0(n24037), .A1(n24036), .B0(n24035), .Y(n25779) );
  INVXL U25356 ( .A(n25674), .Y(n24053) );
  NAND2BX1 U25357 ( .AN(n24040), .B(n6107), .Y(n24041) );
  BUFX3 U25358 ( .A(n24117), .Y(n25761) );
  INVXL U25359 ( .A(n25635), .Y(n24255) );
  AOI211XL U25360 ( .A0(n25761), .A1(n24057), .B0(n24056), .C0(n24055), .Y(
        n2299) );
  AOI21XL U25361 ( .A0(n24374), .A1(n3216), .B0(n24062), .Y(n2114) );
  OAI211X4 U25362 ( .A0(n24067), .A1(n24066), .B0(n24071), .C0(n24065), .Y(
        n24439) );
  INVXL U25363 ( .A(n24070), .Y(n24069) );
  AOI22XL U25364 ( .A0(n24436), .A1(n24073), .B0(n24434), .B1(n24072), .Y(
        n24074) );
  OAI21XL U25365 ( .A0(n24414), .A1(n4572), .B0(n24076), .Y(n2113) );
  AOI222XL U25366 ( .A0(n24417), .A1(n3216), .B0(w1[314]), .B1(n4576), .C0(
        n23088), .C1(w1[346]), .Y(n2112) );
  AOI21XL U25367 ( .A0(n25541), .A1(w1[378]), .B0(n24078), .Y(n1986) );
  OAI21XL U25368 ( .A0(w1[346]), .A1(n25584), .B0(n24079), .Y(n1985) );
  OAI21XL U25369 ( .A0(w1[314]), .A1(n4574), .B0(n24080), .Y(n1984) );
  OAI21XL U25370 ( .A0(n3117), .A1(n26328), .B0(n24081), .Y(n24082) );
  AOI21XL U25371 ( .A0(n25541), .A1(w1[250]), .B0(n24082), .Y(n1858) );
  AOI222XL U25372 ( .A0(n24425), .A1(n25737), .B0(y20[25]), .B1(n25743), .C0(
        n24421), .C1(n20890), .Y(n2385) );
  NAND2XL U25373 ( .A(n24031), .B(n24083), .Y(n24086) );
  ADDHXL U25374 ( .A(n24083), .B(n24304), .CO(n24330), .S(n24084) );
  NAND2XL U25375 ( .A(n25778), .B(n24084), .Y(n24085) );
  NAND3X1 U25376 ( .A(n24086), .B(n24085), .C(n25779), .Y(n25199) );
  AOI21XL U25377 ( .A0(n24048), .A1(n24087), .B0(n3004), .Y(n24088) );
  OAI2BB1X1 U25378 ( .A0N(n3005), .A1N(n24089), .B0(n24088), .Y(n25204) );
  AOI22XL U25379 ( .A0(n24436), .A1(n24093), .B0(n24434), .B1(n24092), .Y(
        n24094) );
  AOI22XL U25380 ( .A0(n25227), .A1(n3025), .B0(y11[24]), .B1(n25025), .Y(
        n24096) );
  AOI21XL U25381 ( .A0(n3060), .A1(n25199), .B0(n24097), .Y(n2480) );
  INVXL U25382 ( .A(n25709), .Y(n24103) );
  OAI21XL U25383 ( .A0(n25120), .A1(n3057), .B0(n24101), .Y(n24102) );
  AOI21XL U25384 ( .A0(n6161), .A1(n24103), .B0(n24102), .Y(n2441) );
  NAND2XL U25385 ( .A(n24031), .B(n24105), .Y(n24108) );
  ADDHXL U25386 ( .A(n24104), .B(n24105), .CO(n25773), .S(n24106) );
  NAND2XL U25387 ( .A(n25778), .B(n24106), .Y(n24107) );
  NAND3X1 U25388 ( .A(n24108), .B(n24107), .C(n25779), .Y(n24396) );
  AOI21XL U25389 ( .A0(n25754), .A1(n24396), .B0(n24113), .Y(n2353) );
  INVXL U25390 ( .A(n24116), .Y(mul5_out[2]) );
  NOR2X1 U25391 ( .A(n24491), .B(n25255), .Y(n24121) );
  INVXL U25392 ( .A(n25590), .Y(n24119) );
  AOI211XL U25393 ( .A0(n3080), .A1(n25591), .B0(n24121), .C0(n24120), .Y(
        n2303) );
  INVXL U25394 ( .A(n24122), .Y(mul5_out[3]) );
  OAI21XL U25395 ( .A0(n3045), .A1(n25907), .B0(n24124), .Y(n24125) );
  AOI211XL U25396 ( .A0(n24127), .A1(n25329), .B0(n24126), .C0(n24125), .Y(
        n2267) );
  AOI21XL U25397 ( .A0(n25754), .A1(n24535), .B0(n24133), .Y(n2307) );
  INVXL U25398 ( .A(n24135), .Y(n24136) );
  OAI21XL U25399 ( .A0(n3045), .A1(n25902), .B0(n24137), .Y(n24138) );
  AOI211XL U25400 ( .A0(n25329), .A1(n24140), .B0(n24139), .C0(n24138), .Y(
        n2269) );
  INVXL U25401 ( .A(n25552), .Y(n24142) );
  AOI211XL U25402 ( .A0(n3080), .A1(n25553), .B0(n24144), .C0(n24143), .Y(
        n2309) );
  AOI21XL U25403 ( .A0(n25754), .A1(n24581), .B0(n24148), .Y(n2311) );
  OAI21XL U25404 ( .A0(n3045), .A1(n25897), .B0(n24150), .Y(n24151) );
  NOR2X1 U25405 ( .A(n24595), .B(n25255), .Y(n24154) );
  AOI211XL U25406 ( .A0(n3080), .A1(n25528), .B0(n24154), .C0(n24153), .Y(
        n2313) );
  INVXL U25407 ( .A(n24155), .Y(n24615) );
  AOI21XL U25408 ( .A0(n25754), .A1(n24615), .B0(n24158), .Y(n2315) );
  OAI21XL U25409 ( .A0(n3045), .A1(n26232), .B0(n24161), .Y(n24162) );
  AOI211XL U25410 ( .A0(n25329), .A1(n24169), .B0(n24163), .C0(n24162), .Y(
        n2273) );
  INVXL U25411 ( .A(n25502), .Y(n24165) );
  AOI211XL U25412 ( .A0(n3080), .A1(n25503), .B0(n24167), .C0(n24166), .Y(
        n2317) );
  INVXL U25413 ( .A(n24169), .Y(n24170) );
  OAI21XL U25414 ( .A0(n3045), .A1(n25905), .B0(n24171), .Y(n24172) );
  AOI211XL U25415 ( .A0(n25329), .A1(n24174), .B0(n24173), .C0(n24172), .Y(
        n2274) );
  AOI21XL U25416 ( .A0(n25754), .A1(n20268), .B0(n24181), .Y(n2321) );
  INVXL U25417 ( .A(n24183), .Y(n24184) );
  OAI21XL U25418 ( .A0(n3045), .A1(n25901), .B0(n24185), .Y(n24186) );
  AOI211XL U25419 ( .A0(n25329), .A1(n24192), .B0(n24187), .C0(n24186), .Y(
        n2276) );
  OAI21XL U25420 ( .A0(n3045), .A1(n26235), .B0(n24193), .Y(n24194) );
  AOI211XL U25421 ( .A0(n25329), .A1(n24201), .B0(n24195), .C0(n24194), .Y(
        n2277) );
  NOR2X1 U25422 ( .A(n24715), .B(n25255), .Y(n24198) );
  AOI211XL U25423 ( .A0(n3080), .A1(n24199), .B0(n24198), .C0(n24197), .Y(
        n2325) );
  INVXL U25424 ( .A(n24200), .Y(mul5_out[14]) );
  INVXL U25425 ( .A(n24201), .Y(n24202) );
  OAI21XL U25426 ( .A0(n3045), .A1(n25899), .B0(n24203), .Y(n24204) );
  AOI211XL U25427 ( .A0(n25329), .A1(n24211), .B0(n24205), .C0(n24204), .Y(
        n2278) );
  NOR2X1 U25428 ( .A(n24744), .B(n25255), .Y(n24209) );
  AOI211XL U25429 ( .A0(n24210), .A1(n3080), .B0(n24209), .C0(n24208), .Y(
        n2327) );
  OAI21XL U25430 ( .A0(n3045), .A1(n25908), .B0(n24212), .Y(n24213) );
  NOR2X1 U25431 ( .A(n24796), .B(n25255), .Y(n24217) );
  OAI21XL U25432 ( .A0(n3045), .A1(n25911), .B0(n24221), .Y(n24222) );
  AOI211XL U25433 ( .A0(n25329), .A1(n24227), .B0(n24223), .C0(n24222), .Y(
        n2280) );
  INVX1 U25434 ( .A(n24224), .Y(n24842) );
  INVXL U25435 ( .A(n24227), .Y(n24228) );
  OAI21XL U25436 ( .A0(n3045), .A1(n25910), .B0(n24229), .Y(n24230) );
  AOI211XL U25437 ( .A0(n25329), .A1(n24237), .B0(n24231), .C0(n24230), .Y(
        n2281) );
  NOR2X1 U25438 ( .A(n24847), .B(n25255), .Y(n24235) );
  OAI21X1 U25439 ( .A0(n24233), .A1(n24256), .B0(n24232), .Y(n24234) );
  AOI211XL U25440 ( .A0(n3080), .A1(n24236), .B0(n24235), .C0(n24234), .Y(
        n2333) );
  OAI21XL U25441 ( .A0(n3045), .A1(n25916), .B0(n24238), .Y(n24239) );
  AOI211XL U25442 ( .A0(n24244), .A1(n3080), .B0(n24243), .C0(n24242), .Y(
        n2335) );
  NOR2X1 U25443 ( .A(n24936), .B(n25255), .Y(n24247) );
  AOI211XL U25444 ( .A0(n25761), .A1(n25379), .B0(n24247), .C0(n24246), .Y(
        n2337) );
  INVXL U25445 ( .A(n24248), .Y(mul5_out[20]) );
  INVXL U25446 ( .A(n24249), .Y(mul5_out[21]) );
  AOI211XL U25447 ( .A0(n25637), .A1(n3080), .B0(n24258), .C0(n24257), .Y(
        n2297) );
  AOI21XL U25448 ( .A0(data[96]), .A1(n4583), .B0(n24266), .Y(n1710) );
  ADDHXL U25449 ( .A(n24268), .B(n24269), .CO(n24382), .S(n24270) );
  NAND2XL U25450 ( .A(n24031), .B(n24280), .Y(n24283) );
  ADDHXL U25451 ( .A(n24279), .B(n24280), .CO(n24104), .S(n24281) );
  NAND2XL U25452 ( .A(n25778), .B(n24281), .Y(n24282) );
  INVXL U25453 ( .A(n25170), .Y(n24290) );
  ADDHXL U25454 ( .A(n24284), .B(n24285), .CO(n24375), .S(n24287) );
  AOI21XL U25455 ( .A0(n24048), .A1(n24285), .B0(n3004), .Y(n24286) );
  OAI2BB1X1 U25456 ( .A0N(n3005), .A1N(n24287), .B0(n24286), .Y(n25174) );
  AOI222XL U25457 ( .A0(n25083), .A1(n25292), .B0(in_valid_w2), .B1(
        weight2[27]), .C0(w2[91]), .C1(n25822), .Y(n2227) );
  AOI22XL U25458 ( .A0(n24436), .A1(n24296), .B0(n24434), .B1(n24295), .Y(
        n24297) );
  AOI222XL U25459 ( .A0(n25090), .A1(n25292), .B0(w2[59]), .B1(n25822), .C0(
        w2[91]), .C1(in_valid_w2), .Y(n2195) );
  AOI22XL U25460 ( .A0(n24436), .A1(n24301), .B0(n24434), .B1(n24300), .Y(
        n24302) );
  AOI222XL U25461 ( .A0(n25816), .A1(n25292), .B0(w2[62]), .B1(n25822), .C0(
        w2[94]), .C1(in_valid_w2), .Y(n2198) );
  NAND2XL U25462 ( .A(n24031), .B(n24304), .Y(n24307) );
  NAND2XL U25463 ( .A(n25778), .B(n24305), .Y(n24306) );
  AOI22XL U25464 ( .A0(n24436), .A1(n24310), .B0(n24434), .B1(n24309), .Y(
        n24311) );
  AOI22XL U25465 ( .A0(n25810), .A1(n3025), .B0(y11[23]), .B1(n24739), .Y(
        n24313) );
  AOI21XL U25466 ( .A0(n3060), .A1(n25803), .B0(n24314), .Y(n2479) );
  OAI21XL U25467 ( .A0(n24317), .A1(n3057), .B0(n24316), .Y(n24318) );
  AOI21XL U25468 ( .A0(n24525), .A1(n24319), .B0(n24318), .Y(n2439) );
  OAI21XL U25469 ( .A0(n25810), .A1(n4571), .B0(n24320), .Y(n2101) );
  AOI222XL U25470 ( .A0(n24321), .A1(n3216), .B0(w1[311]), .B1(n4578), .C0(
        n3061), .C1(w1[343]), .Y(n2100) );
  OAI21XL U25471 ( .A0(w1[343]), .A1(n3226), .B0(n24322), .Y(n1973) );
  AOI21XL U25472 ( .A0(n24325), .A1(n3216), .B0(n24324), .Y(n2102) );
  AOI21XL U25473 ( .A0(n25541), .A1(w1[375]), .B0(n24327), .Y(n1974) );
  OAI21XL U25474 ( .A0(n3117), .A1(n26329), .B0(n24328), .Y(n24329) );
  AOI21XL U25475 ( .A0(n25541), .A1(w1[247]), .B0(n24329), .Y(n1846) );
  NAND2XL U25476 ( .A(n24031), .B(n24331), .Y(n24334) );
  ADDHXL U25477 ( .A(n24330), .B(n24331), .CO(n24409), .S(n24332) );
  NAND2XL U25478 ( .A(n25778), .B(n24332), .Y(n24333) );
  NAND3X1 U25479 ( .A(n24334), .B(n24333), .C(n25779), .Y(n25191) );
  AOI21XL U25480 ( .A0(n24048), .A1(n24336), .B0(n3004), .Y(n24337) );
  OAI2BB1X1 U25481 ( .A0N(n3005), .A1N(n24338), .B0(n24337), .Y(n25195) );
  AOI22XL U25482 ( .A0(n24436), .A1(n24342), .B0(n24434), .B1(n24341), .Y(
        n24343) );
  AOI22XL U25483 ( .A0(n24373), .A1(n3025), .B0(y11[25]), .B1(n25025), .Y(
        n24345) );
  AOI21XL U25484 ( .A0(n25675), .A1(n25191), .B0(n24346), .Y(n2481) );
  INVXL U25485 ( .A(n24352), .Y(n24358) );
  OAI21XL U25486 ( .A0(n24363), .A1(n3057), .B0(n24356), .Y(n24357) );
  AOI21XL U25487 ( .A0(n6161), .A1(n24358), .B0(n24357), .Y(n2443) );
  AOI21XL U25488 ( .A0(n25220), .A1(n24361), .B0(n25219), .Y(n24362) );
  OAI2BB1X1 U25489 ( .A0N(n25099), .A1N(n23643), .B0(n24362), .Y(mul5_out[25])
         );
  INVXL U25490 ( .A(n24363), .Y(n24370) );
  AOI222XL U25491 ( .A0(n24370), .A1(n25292), .B0(in_valid_w2), .B1(
        weight2[25]), .C0(w2[89]), .C1(n25822), .Y(n2225) );
  AOI21XL U25492 ( .A0(n25541), .A1(w1[377]), .B0(n24365), .Y(n1982) );
  OAI21XL U25493 ( .A0(n3117), .A1(n26330), .B0(n24366), .Y(n24367) );
  AOI21XL U25494 ( .A0(n25541), .A1(w1[249]), .B0(n24367), .Y(n1854) );
  AOI21XL U25495 ( .A0(n24370), .A1(n3216), .B0(n24369), .Y(n2110) );
  OAI21XL U25496 ( .A0(n24373), .A1(n4574), .B0(n24371), .Y(n2109) );
  OAI21XL U25497 ( .A0(w1[345]), .A1(n4571), .B0(n24372), .Y(n1981) );
  AOI222XL U25498 ( .A0(n24373), .A1(n25292), .B0(w2[57]), .B1(n25822), .C0(
        w2[89]), .C1(in_valid_w2), .Y(n2193) );
  AOI222XL U25499 ( .A0(n24374), .A1(n25292), .B0(in_valid_w2), .B1(
        weight2[26]), .C0(w2[90]), .C1(n25822), .Y(n2226) );
  AOI222XL U25500 ( .A0(n24414), .A1(n25292), .B0(w2[58]), .B1(n25822), .C0(
        w2[90]), .C1(in_valid_w2), .Y(n2194) );
  ADDHXL U25501 ( .A(n24375), .B(n24376), .CO(n25788), .S(n24378) );
  AOI21XL U25502 ( .A0(n24048), .A1(n24376), .B0(n3004), .Y(n24377) );
  OAI2BB1X1 U25503 ( .A0N(n3005), .A1N(n24378), .B0(n24377), .Y(n25166) );
  ADDHXL U25504 ( .A(n24382), .B(n24383), .CO(n23660), .S(n24384) );
  AOI22XL U25505 ( .A0(n24436), .A1(n24391), .B0(n24434), .B1(n24390), .Y(
        n24392) );
  AOI22XL U25506 ( .A0(n24459), .A1(n3025), .B0(y11[28]), .B1(n24739), .Y(
        n24394) );
  AOI21XL U25507 ( .A0(n3060), .A1(n24396), .B0(n24395), .Y(n2484) );
  INVXL U25508 ( .A(n24449), .Y(n24404) );
  OAI21XL U25509 ( .A0(n24405), .A1(n3057), .B0(n24402), .Y(n24403) );
  AOI21XL U25510 ( .A0(n3060), .A1(n24404), .B0(n24403), .Y(n2449) );
  AOI222XL U25511 ( .A0(n24456), .A1(n25292), .B0(in_valid_w2), .B1(
        weight2[28]), .C0(w2[92]), .C1(n25822), .Y(n2228) );
  INVXL U25512 ( .A(n25080), .Y(n24407) );
  AOI21XL U25513 ( .A0(n25076), .A1(n24525), .B0(n24408), .Y(n2446) );
  NAND2XL U25514 ( .A(n24031), .B(n24410), .Y(n24413) );
  ADDHXL U25515 ( .A(n24409), .B(n24410), .CO(n24279), .S(n24411) );
  NAND2XL U25516 ( .A(n25778), .B(n24411), .Y(n24412) );
  AOI22XL U25517 ( .A0(n24414), .A1(n3025), .B0(y11[26]), .B1(n24958), .Y(
        n24415) );
  AOI21XL U25518 ( .A0(n3060), .A1(n25678), .B0(n24416), .Y(n2482) );
  INVXL U25519 ( .A(n24417), .Y(n24419) );
  AOI21XL U25520 ( .A0(n25720), .A1(n24525), .B0(n24420), .Y(n2444) );
  INVXL U25521 ( .A(n24421), .Y(n24423) );
  AOI21XL U25522 ( .A0(n24425), .A1(n24525), .B0(n24424), .Y(n2442) );
  AOI222XL U25523 ( .A0(n25113), .A1(n25292), .B0(in_valid_w2), .B1(
        weight2[29]), .C0(w2[93]), .C1(n25822), .Y(n2229) );
  AOI22XL U25524 ( .A0(n24436), .A1(n24435), .B0(n24434), .B1(n24433), .Y(
        n24437) );
  AOI222XL U25525 ( .A0(n25671), .A1(n25292), .B0(w2[61]), .B1(n25822), .C0(
        w2[93]), .C1(in_valid_w2), .Y(n2197) );
  OAI21XL U25526 ( .A0(n25832), .A1(n24440), .B0(n25829), .Y(n24444) );
  INVXL U25527 ( .A(n24440), .Y(n24441) );
  NOR3XL U25528 ( .A(n25832), .B(n24443), .C(n24441), .Y(n24442) );
  AOI21XL U25529 ( .A0(n24447), .A1(in_valid_d), .B0(n24446), .Y(n24448) );
  OAI21XL U25530 ( .A0(n3117), .A1(n26331), .B0(n24452), .Y(n24453) );
  AOI21XL U25531 ( .A0(n25541), .A1(w1[252]), .B0(n24453), .Y(n1866) );
  AOI21XL U25532 ( .A0(n24456), .A1(n3216), .B0(n24455), .Y(n2122) );
  OAI21XL U25533 ( .A0(n24459), .A1(n3226), .B0(n24457), .Y(n2121) );
  OAI21XL U25534 ( .A0(w1[348]), .A1(n25584), .B0(n24458), .Y(n1993) );
  AOI222XL U25535 ( .A0(n24459), .A1(n25292), .B0(w2[60]), .B1(n25822), .C0(
        w2[92]), .C1(in_valid_w2), .Y(n2196) );
  CLKINVX3 U25536 ( .A(n25693), .Y(n25675) );
  INVXL U25537 ( .A(n24460), .Y(n24466) );
  INVXL U25538 ( .A(n24462), .Y(n24461) );
  AOI22XL U25539 ( .A0(n25677), .A1(n25664), .B0(n24958), .B1(y11[0]), .Y(
        n24464) );
  AOI21XL U25540 ( .A0(n25675), .A1(n24466), .B0(n24465), .Y(n2456) );
  XNOR2XL U25541 ( .A(n24467), .B(n25138), .Y(n24468) );
  OAI21XL U25542 ( .A0(n25625), .A1(n3227), .B0(n24470), .Y(n24471) );
  OAI21XL U25543 ( .A0(n24473), .A1(n3227), .B0(n24472), .Y(n24474) );
  AOI21XL U25544 ( .A0(n24475), .A1(n24525), .B0(n24474), .Y(n2394) );
  AOI22XL U25545 ( .A0(n25609), .A1(n3025), .B0(n24739), .B1(y11[2]), .Y(
        n24480) );
  OAI21XL U25546 ( .A0(n25611), .A1(n3057), .B0(n24485), .Y(n24486) );
  OAI21XL U25547 ( .A0(n24488), .A1(n3057), .B0(n24487), .Y(n24489) );
  AOI21XL U25548 ( .A0(n24490), .A1(n24525), .B0(n24489), .Y(n2396) );
  INVXL U25549 ( .A(n24491), .Y(n24501) );
  AOI22XL U25550 ( .A0(n25596), .A1(n3025), .B0(n24958), .B1(y11[3]), .Y(
        n24499) );
  AOI21XL U25551 ( .A0(n25675), .A1(n24501), .B0(n24500), .Y(n2459) );
  INVXL U25552 ( .A(n25594), .Y(n24510) );
  INVXL U25553 ( .A(n24507), .Y(n24504) );
  OAI21XL U25554 ( .A0(n25598), .A1(n3057), .B0(n24508), .Y(n24509) );
  OAI21XL U25555 ( .A0(n24512), .A1(n3057), .B0(n24511), .Y(n24513) );
  AOI21XL U25556 ( .A0(n24514), .A1(n24525), .B0(n24513), .Y(n2398) );
  INVXL U25557 ( .A(n24515), .Y(n24521) );
  OAI21XL U25558 ( .A0(n25579), .A1(n3057), .B0(n24519), .Y(n24520) );
  AOI21XL U25559 ( .A0(n24521), .A1(n24525), .B0(n24520), .Y(n2401) );
  OAI21XL U25560 ( .A0(n24523), .A1(n3057), .B0(n24522), .Y(n24524) );
  AOI21XL U25561 ( .A0(n24526), .A1(n24525), .B0(n24524), .Y(n2400) );
  NOR2XL U25562 ( .A(n24572), .B(n24527), .Y(n24529) );
  INVXL U25563 ( .A(n24531), .Y(n24528) );
  AOI22XL U25564 ( .A0(n25566), .A1(n25664), .B0(n24958), .B1(y11[5]), .Y(
        n24533) );
  AOI21XL U25565 ( .A0(n25675), .A1(n24535), .B0(n24534), .Y(n2461) );
  INVXL U25566 ( .A(n24536), .Y(n24544) );
  INVXL U25567 ( .A(n24541), .Y(n24538) );
  OAI21XL U25568 ( .A0(n25569), .A1(n3057), .B0(n24542), .Y(n24543) );
  AOI21XL U25569 ( .A0(n24544), .A1(n25675), .B0(n24543), .Y(n2403) );
  OAI21XL U25570 ( .A0(n24546), .A1(n3057), .B0(n24545), .Y(n24547) );
  NOR2XL U25571 ( .A(n24572), .B(n24569), .Y(n24550) );
  INVXL U25572 ( .A(n24570), .Y(n24549) );
  AOI22XL U25573 ( .A0(n25558), .A1(n25664), .B0(n24958), .B1(y11[6]), .Y(
        n24553) );
  AOI21XL U25574 ( .A0(n25675), .A1(n24555), .B0(n24554), .Y(n2462) );
  NOR2XL U25575 ( .A(n24586), .B(n24583), .Y(n24557) );
  AOI22X1 U25576 ( .A0(n3029), .A1(n24584), .B0(n25290), .B1(n24558), .Y(
        n25559) );
  OAI21XL U25577 ( .A0(n25559), .A1(n3057), .B0(n24559), .Y(n24560) );
  AOI21XL U25578 ( .A0(n11478), .A1(n25675), .B0(n24560), .Y(n2405) );
  NOR2XL U25579 ( .A(n24562), .B(n24561), .Y(n24564) );
  INVXL U25580 ( .A(n24566), .Y(n24563) );
  XNOR2X1 U25581 ( .A(n24564), .B(n24563), .Y(n24565) );
  OAI21XL U25582 ( .A0(n25308), .A1(n3057), .B0(n24567), .Y(n24568) );
  AOI21XL U25583 ( .A0(n25740), .A1(n25675), .B0(n24568), .Y(n2404) );
  INVXL U25584 ( .A(n24569), .Y(n24571) );
  NAND2XL U25585 ( .A(n24571), .B(n24570), .Y(n24573) );
  NOR2XL U25586 ( .A(n24573), .B(n24572), .Y(n24575) );
  AOI22XL U25587 ( .A0(n25545), .A1(n3025), .B0(n24958), .B1(y11[7]), .Y(
        n24579) );
  OAI21X1 U25588 ( .A0(n24582), .A1(n3059), .B0(n24579), .Y(n24580) );
  AOI21XL U25589 ( .A0(n3060), .A1(n24581), .B0(n24580), .Y(n2463) );
  INVXL U25590 ( .A(n24582), .Y(n24594) );
  AOI22X1 U25591 ( .A0(n3029), .A1(n24591), .B0(n25290), .B1(n24590), .Y(
        n25547) );
  OAI21XL U25592 ( .A0(n25547), .A1(n3057), .B0(n24592), .Y(n24593) );
  AOI21XL U25593 ( .A0(n24594), .A1(n3060), .B0(n24593), .Y(n2407) );
  INVXL U25594 ( .A(n24595), .Y(n24601) );
  AOI21XL U25595 ( .A0(n25675), .A1(n24601), .B0(n24600), .Y(n2464) );
  XNOR2X1 U25596 ( .A(n24775), .B(n24602), .Y(n24603) );
  OAI21XL U25597 ( .A0(n25536), .A1(n3057), .B0(n24604), .Y(n24605) );
  NAND2XL U25598 ( .A(n24760), .B(n24607), .Y(n24609) );
  AOI22XL U25599 ( .A0(n25518), .A1(n25664), .B0(n24958), .B1(y11[9]), .Y(
        n24613) );
  AOI21XL U25600 ( .A0(n3060), .A1(n24615), .B0(n24614), .Y(n2465) );
  INVXL U25601 ( .A(n24616), .Y(n24625) );
  NAND2XL U25602 ( .A(n24775), .B(n24618), .Y(n24620) );
  OAI21XL U25603 ( .A0(n25521), .A1(n3057), .B0(n24623), .Y(n24624) );
  AOI21XL U25604 ( .A0(n24625), .A1(n25675), .B0(n24624), .Y(n2411) );
  INVX1 U25605 ( .A(n24626), .Y(n24633) );
  NAND2XL U25606 ( .A(n24760), .B(n24627), .Y(n24628) );
  INVXL U25607 ( .A(n25506), .Y(n24640) );
  NAND2XL U25608 ( .A(n24775), .B(n24634), .Y(n24635) );
  OAI21XL U25609 ( .A0(n25510), .A1(n3057), .B0(n24638), .Y(n24639) );
  AOI21XL U25610 ( .A0(n24640), .A1(n3060), .B0(n24639), .Y(n2413) );
  OAI21XL U25611 ( .A0(n24642), .A1(n3057), .B0(n24641), .Y(n24643) );
  AOI21XL U25612 ( .A0(n24644), .A1(n24525), .B0(n24643), .Y(n2412) );
  NAND2XL U25613 ( .A(n24760), .B(n24647), .Y(n24649) );
  AOI22XL U25614 ( .A0(n25495), .A1(n25664), .B0(n24958), .B1(y11[11]), .Y(
        n24653) );
  AOI21XL U25615 ( .A0(n25675), .A1(n24655), .B0(n24654), .Y(n2467) );
  INVXL U25616 ( .A(n24656), .Y(n24666) );
  NAND2XL U25617 ( .A(n24775), .B(n24659), .Y(n24661) );
  XOR2X1 U25618 ( .A(n24661), .B(n24660), .Y(n24662) );
  AOI22XL U25619 ( .A0(n24739), .A1(y12[11]), .B0(n3120), .B1(y11[11]), .Y(
        n24664) );
  OAI21XL U25620 ( .A0(n25497), .A1(n3057), .B0(n24664), .Y(n24665) );
  AOI21XL U25621 ( .A0(n24666), .A1(n25675), .B0(n24665), .Y(n2415) );
  NAND2XL U25622 ( .A(n24775), .B(n24667), .Y(n24668) );
  XOR2X1 U25623 ( .A(n24668), .B(n24698), .Y(n24669) );
  OAI21XL U25624 ( .A0(n25487), .A1(n3057), .B0(n24671), .Y(n24672) );
  AOI21XL U25625 ( .A0(n24673), .A1(n3060), .B0(n24672), .Y(n2417) );
  AOI22XL U25626 ( .A0(n24739), .A1(y10[12]), .B0(n3120), .B1(y12[12]), .Y(
        n24674) );
  OAI21XL U25627 ( .A0(n24675), .A1(n3057), .B0(n24674), .Y(n24676) );
  NOR2XL U25628 ( .A(n3030), .B(n24678), .Y(n24679) );
  AOI21XL U25629 ( .A0(n24680), .A1(n3030), .B0(n24679), .Y(n24749) );
  NOR2XL U25630 ( .A(n24681), .B(n3032), .Y(n24682) );
  AOI21XL U25631 ( .A0(n24749), .A1(n3032), .B0(n24682), .Y(n24825) );
  NAND2XL U25632 ( .A(n24994), .B(n3075), .Y(n24686) );
  INVXL U25633 ( .A(n24811), .Y(n24758) );
  NOR2XL U25634 ( .A(n24758), .B(n24688), .Y(n24689) );
  NAND2XL U25635 ( .A(n24689), .B(n24760), .Y(n24690) );
  AOI22XL U25636 ( .A0(n25472), .A1(n25664), .B0(n24958), .B1(y11[13]), .Y(
        n24694) );
  AOI21XL U25637 ( .A0(n3060), .A1(n24696), .B0(n24695), .Y(n2469) );
  NOR2XL U25638 ( .A(n24773), .B(n24698), .Y(n24699) );
  NAND2XL U25639 ( .A(n24699), .B(n24775), .Y(n24701) );
  OAI21XL U25640 ( .A0(n25473), .A1(n3057), .B0(n24704), .Y(n24705) );
  AOI21XL U25641 ( .A0(n24706), .A1(n3060), .B0(n24705), .Y(n2419) );
  NOR2XL U25642 ( .A(n24787), .B(n24707), .Y(n24708) );
  NAND2XL U25643 ( .A(n24708), .B(n24789), .Y(n24710) );
  OAI21XL U25644 ( .A0(n25316), .A1(n3057), .B0(n24713), .Y(n24714) );
  AOI21XL U25645 ( .A0(n25738), .A1(n3060), .B0(n24714), .Y(n2418) );
  INVXL U25646 ( .A(n24715), .Y(n24734) );
  NAND2XL U25647 ( .A(n3030), .B(n24717), .Y(n24718) );
  OAI21XL U25648 ( .A0(n3030), .A1(n24746), .B0(n24718), .Y(n24800) );
  OAI22XL U25649 ( .A0(n3072), .A1(n24800), .B0(n24719), .B1(n20138), .Y(
        n24853) );
  OAI22XL U25650 ( .A0(n20182), .A1(n24853), .B0(n24720), .B1(n3069), .Y(
        n25340) );
  NOR2XL U25651 ( .A(n25340), .B(n20066), .Y(n24724) );
  NOR2XL U25652 ( .A(n24721), .B(n3075), .Y(n24723) );
  NAND2XL U25653 ( .A(n24726), .B(n24725), .Y(n24809) );
  NOR2XL U25654 ( .A(n24758), .B(n24809), .Y(n24727) );
  NAND2XL U25655 ( .A(n24727), .B(n24760), .Y(n24729) );
  XOR2X1 U25656 ( .A(n24729), .B(n24728), .Y(n24730) );
  INVX1 U25657 ( .A(n24731), .Y(n25459) );
  AOI22XL U25658 ( .A0(n25459), .A1(n3025), .B0(n24958), .B1(y11[14]), .Y(
        n24732) );
  OAI21X1 U25659 ( .A0(n24735), .A1(n3024), .B0(n24732), .Y(n24733) );
  AOI21XL U25660 ( .A0(n24525), .A1(n24734), .B0(n24733), .Y(n2470) );
  OAI21XL U25661 ( .A0(n25461), .A1(n3057), .B0(n24736), .Y(n24737) );
  AOI22XL U25662 ( .A0(n24739), .A1(y10[14]), .B0(n3120), .B1(y12[14]), .Y(
        n24740) );
  OAI21XL U25663 ( .A0(n24741), .A1(n3057), .B0(n24740), .Y(n24742) );
  INVXL U25664 ( .A(n24744), .Y(n24768) );
  NOR2XL U25665 ( .A(n3030), .B(n24745), .Y(n24748) );
  NOR2XL U25666 ( .A(n24748), .B(n24747), .Y(n24829) );
  AOI22XL U25667 ( .A0(n24749), .A1(n3072), .B0(n24829), .B1(n20138), .Y(
        n24895) );
  NAND2XL U25668 ( .A(n3069), .B(n24895), .Y(n24750) );
  OAI21XL U25669 ( .A0(n3069), .A1(n24751), .B0(n24750), .Y(n24754) );
  NAND2XL U25670 ( .A(n24752), .B(n20066), .Y(n24753) );
  OAI21XL U25671 ( .A0(n3074), .A1(n24756), .B0(n24755), .Y(n24807) );
  INVXL U25672 ( .A(n24809), .Y(n24757) );
  NAND2XL U25673 ( .A(n24757), .B(n24808), .Y(n24759) );
  NOR2XL U25674 ( .A(n24759), .B(n24758), .Y(n24761) );
  NAND2XL U25675 ( .A(n24761), .B(n24760), .Y(n24763) );
  AOI22XL U25676 ( .A0(n25448), .A1(n3025), .B0(n24958), .B1(y11[15]), .Y(
        n24766) );
  AOI21XL U25677 ( .A0(n3060), .A1(n24768), .B0(n24767), .Y(n2471) );
  INVXL U25678 ( .A(n24770), .Y(n24772) );
  NAND2XL U25679 ( .A(n24772), .B(n24771), .Y(n24774) );
  NOR2XL U25680 ( .A(n24774), .B(n24773), .Y(n24776) );
  NAND2XL U25681 ( .A(n24776), .B(n24775), .Y(n24778) );
  AOI22XL U25682 ( .A0(n25025), .A1(y12[15]), .B0(n3120), .B1(y11[15]), .Y(
        n24781) );
  OAI21XL U25683 ( .A0(n25449), .A1(n3057), .B0(n24781), .Y(n24782) );
  AOI21XL U25684 ( .A0(n20776), .A1(n3060), .B0(n24782), .Y(n2423) );
  NOR2XL U25685 ( .A(n24788), .B(n24787), .Y(n24790) );
  NAND2XL U25686 ( .A(n24790), .B(n24789), .Y(n24791) );
  OAI21XL U25687 ( .A0(n25319), .A1(n3057), .B0(n24794), .Y(n24795) );
  AOI21XL U25688 ( .A0(n25735), .A1(n3060), .B0(n24795), .Y(n2422) );
  INVXL U25689 ( .A(n24796), .Y(n24820) );
  NOR2XL U25690 ( .A(n24797), .B(n3075), .Y(n24806) );
  NAND2XL U25691 ( .A(n3030), .B(n24798), .Y(n24799) );
  OAI21XL U25692 ( .A0(n3030), .A1(n20096), .B0(n24799), .Y(n24852) );
  OAI22XL U25693 ( .A0(n3072), .A1(n24852), .B0(n24800), .B1(n20138), .Y(
        n24943) );
  OAI21XL U25694 ( .A0(n24943), .A1(n20182), .B0(n3075), .Y(n24803) );
  NOR2XL U25695 ( .A(n24801), .B(n3069), .Y(n24802) );
  NAND2XL U25696 ( .A(n24808), .B(n24807), .Y(n24810) );
  NOR2XL U25697 ( .A(n24810), .B(n24809), .Y(n24812) );
  NOR2X2 U25698 ( .A(n24814), .B(n24813), .Y(n25358) );
  AOI22XL U25699 ( .A0(n25435), .A1(n3025), .B0(n25025), .B1(y11[16]), .Y(
        n24818) );
  AOI21XL U25700 ( .A0(n3060), .A1(n24820), .B0(n24819), .Y(n2472) );
  INVXL U25701 ( .A(n24821), .Y(n24824) );
  OAI21XL U25702 ( .A0(n25437), .A1(n3057), .B0(n24822), .Y(n24823) );
  NAND2XL U25703 ( .A(n24825), .B(n24894), .Y(n24831) );
  NOR2XL U25704 ( .A(n3030), .B(n24826), .Y(n24827) );
  AOI21XL U25705 ( .A0(n24828), .A1(n3030), .B0(n24827), .Y(n24893) );
  AOI22XL U25706 ( .A0(n24893), .A1(n3032), .B0(n24829), .B1(n3072), .Y(n24993) );
  AOI21XL U25707 ( .A0(n24993), .A1(n3069), .B0(n20066), .Y(n24830) );
  OAI21XL U25708 ( .A0(n3075), .A1(n24833), .B0(n24832), .Y(n24834) );
  OAI21XL U25709 ( .A0(n24835), .A1(n3074), .B0(n24834), .Y(n24859) );
  NAND2XL U25710 ( .A(n25358), .B(n24860), .Y(n24837) );
  XOR2X1 U25711 ( .A(n24837), .B(n24836), .Y(n24838) );
  AOI22XL U25712 ( .A0(n25421), .A1(n25664), .B0(n24958), .B1(y11[17]), .Y(
        n24840) );
  AOI21XL U25713 ( .A0(n24525), .A1(n24842), .B0(n24841), .Y(n2473) );
  INVXL U25714 ( .A(n24843), .Y(n24846) );
  OAI21XL U25715 ( .A0(n25423), .A1(n3057), .B0(n24844), .Y(n24845) );
  AOI21XL U25716 ( .A0(n24846), .A1(n6161), .B0(n24845), .Y(n2427) );
  NOR2XL U25717 ( .A(n24848), .B(n3075), .Y(n24858) );
  NAND2XL U25718 ( .A(n3030), .B(n24849), .Y(n24850) );
  OAI21XL U25719 ( .A0(n3030), .A1(n24851), .B0(n24850), .Y(n24940) );
  OAI22XL U25720 ( .A0(n3072), .A1(n24940), .B0(n24852), .B1(n20138), .Y(
        n25341) );
  OAI21XL U25721 ( .A0(n25341), .A1(n20182), .B0(n3075), .Y(n24855) );
  NOR2XL U25722 ( .A(n24853), .B(n3069), .Y(n24854) );
  NAND2XL U25723 ( .A(n24860), .B(n24859), .Y(n24953) );
  NAND2XL U25724 ( .A(n25358), .B(n24861), .Y(n24862) );
  XOR2X1 U25725 ( .A(n24862), .B(n24903), .Y(n24863) );
  AOI22XL U25726 ( .A0(n25407), .A1(n25664), .B0(n24958), .B1(y11[18]), .Y(
        n24865) );
  AOI21XL U25727 ( .A0(n3060), .A1(n24867), .B0(n24866), .Y(n2474) );
  INVXL U25728 ( .A(n24868), .Y(n24887) );
  NAND2XL U25729 ( .A(n25271), .B(n24871), .Y(n24872) );
  OAI21XL U25730 ( .A0(n25269), .A1(n15716), .B0(n24872), .Y(n24964) );
  OAI22XL U25731 ( .A0(n3127), .A1(n24964), .B0(n24873), .B1(n25273), .Y(
        n25266) );
  OAI21XL U25732 ( .A0(n25266), .A1(n15808), .B0(n3077), .Y(n24876) );
  NOR2XL U25733 ( .A(n24874), .B(n3125), .Y(n24875) );
  NAND2XL U25734 ( .A(n4782), .B(n24880), .Y(n24977) );
  NAND2XL U25735 ( .A(n25286), .B(n24882), .Y(n24883) );
  OAI21XL U25736 ( .A0(n25408), .A1(n3057), .B0(n24885), .Y(n24886) );
  OAI21XL U25737 ( .A0(n3030), .A1(n24891), .B0(n24890), .Y(n24989) );
  OAI21XL U25738 ( .A0(n24989), .A1(n3072), .B0(n3069), .Y(n24892) );
  NAND2XL U25739 ( .A(n24898), .B(n20066), .Y(n24899) );
  OAI21XL U25740 ( .A0(n24902), .A1(n3074), .B0(n24901), .Y(n24950) );
  NOR2XL U25741 ( .A(n24953), .B(n24903), .Y(n24904) );
  NAND2XL U25742 ( .A(n25358), .B(n24904), .Y(n24906) );
  XOR2X1 U25743 ( .A(n24906), .B(n24905), .Y(n24907) );
  AOI22XL U25744 ( .A0(n25392), .A1(n25664), .B0(n24739), .B1(y11[19]), .Y(
        n24910) );
  OAI21X1 U25745 ( .A0(n24913), .A1(n3024), .B0(n24910), .Y(n24911) );
  AOI21XL U25746 ( .A0(n24525), .A1(n24912), .B0(n24911), .Y(n2475) );
  INVXL U25747 ( .A(n24913), .Y(n24935) );
  NAND2XL U25748 ( .A(n24914), .B(n15808), .Y(n24923) );
  NOR2XL U25749 ( .A(n25269), .B(n3133), .Y(n24916) );
  AOI21XL U25750 ( .A0(n25011), .A1(n3070), .B0(n24917), .Y(n24921) );
  OAI21XL U25751 ( .A0(n24925), .A1(n3077), .B0(n24924), .Y(n24926) );
  OAI21XL U25752 ( .A0(n24927), .A1(n3076), .B0(n24926), .Y(n24974) );
  NOR2XL U25753 ( .A(n24977), .B(n24928), .Y(n24929) );
  NAND2XL U25754 ( .A(n25286), .B(n24929), .Y(n24931) );
  XOR2X1 U25755 ( .A(n24931), .B(n24930), .Y(n24932) );
  OAI21XL U25756 ( .A0(n25394), .A1(n3057), .B0(n24933), .Y(n24934) );
  AOI21XL U25757 ( .A0(n24935), .A1(n6161), .B0(n24934), .Y(n2431) );
  INVXL U25758 ( .A(n24936), .Y(n24961) );
  NAND2XL U25759 ( .A(n3030), .B(n24938), .Y(n24939) );
  OAI21XL U25760 ( .A0(n3030), .A1(n20100), .B0(n24939), .Y(n25342) );
  NOR2XL U25761 ( .A(n25342), .B(n3072), .Y(n24942) );
  NOR2XL U25762 ( .A(n24940), .B(n20138), .Y(n24941) );
  OAI21XL U25763 ( .A0(n24942), .A1(n24941), .B0(n3075), .Y(n24945) );
  NOR2XL U25764 ( .A(n24943), .B(n3069), .Y(n24944) );
  OAI21XL U25765 ( .A0(n24947), .A1(n3075), .B0(n24946), .Y(n24948) );
  OAI21XL U25766 ( .A0(n24949), .A1(n3074), .B0(n24948), .Y(n24956) );
  NAND2XL U25767 ( .A(n24951), .B(n24950), .Y(n24952) );
  NAND2XL U25768 ( .A(n25358), .B(n25356), .Y(n24954) );
  AOI22XL U25769 ( .A0(n25384), .A1(n25664), .B0(n24958), .B1(y11[20]), .Y(
        n24959) );
  OAI21X1 U25770 ( .A0(n25382), .A1(n3024), .B0(n24959), .Y(n24960) );
  AOI21XL U25771 ( .A0(n24525), .A1(n24961), .B0(n24960), .Y(n2476) );
  INVXL U25772 ( .A(n25382), .Y(n24983) );
  NAND2XL U25773 ( .A(n25271), .B(n24962), .Y(n24963) );
  OAI21XL U25774 ( .A0(n25271), .A1(n3135), .B0(n24963), .Y(n25267) );
  NOR2XL U25775 ( .A(n24964), .B(n3070), .Y(n24965) );
  OAI21XL U25776 ( .A0(n24966), .A1(n24965), .B0(n3077), .Y(n24969) );
  NOR2XL U25777 ( .A(n24967), .B(n3125), .Y(n24968) );
  OAI21XL U25778 ( .A0(n24971), .A1(n3077), .B0(n24970), .Y(n24972) );
  OAI21XL U25779 ( .A0(n24973), .A1(n3076), .B0(n24972), .Y(n24980) );
  NAND2XL U25780 ( .A(n24975), .B(n24974), .Y(n24976) );
  NAND2XL U25781 ( .A(n25286), .B(n25284), .Y(n24978) );
  OAI21XL U25782 ( .A0(n25386), .A1(n3057), .B0(n24981), .Y(n24982) );
  OAI21XL U25783 ( .A0(n24991), .A1(n24990), .B0(n3075), .Y(n24992) );
  NAND2XL U25784 ( .A(n24994), .B(n20066), .Y(n24995) );
  OAI21XL U25785 ( .A0(n24998), .A1(n3074), .B0(n24997), .Y(n25003) );
  INVXL U25786 ( .A(n25356), .Y(n24999) );
  NOR2XL U25787 ( .A(n24999), .B(n25353), .Y(n25000) );
  NAND2XL U25788 ( .A(n25358), .B(n25000), .Y(n25001) );
  INVXL U25789 ( .A(n25003), .Y(n25354) );
  XOR2X1 U25790 ( .A(n25001), .B(n25354), .Y(n25002) );
  AOI22XL U25791 ( .A0(n25371), .A1(n25664), .B0(n24958), .B1(y11[21]), .Y(
        n25005) );
  INVXL U25792 ( .A(n25731), .Y(n25028) );
  NOR2XL U25793 ( .A(n25006), .B(n3077), .Y(n25018) );
  OAI21XL U25794 ( .A0(n25015), .A1(n3125), .B0(n25014), .Y(n25016) );
  INVXL U25795 ( .A(n25016), .Y(n25017) );
  OAI22XL U25796 ( .A0(n25019), .A1(n3076), .B0(n25018), .B1(n25017), .Y(
        n25024) );
  INVXL U25797 ( .A(n25284), .Y(n25020) );
  NOR2XL U25798 ( .A(n25020), .B(n25281), .Y(n25021) );
  NAND2XL U25799 ( .A(n25286), .B(n25021), .Y(n25022) );
  INVXL U25800 ( .A(n25024), .Y(n25282) );
  XOR2X1 U25801 ( .A(n25022), .B(n25282), .Y(n25023) );
  OAI21XL U25802 ( .A0(n25373), .A1(n3057), .B0(n25026), .Y(n25027) );
  AOI21XL U25803 ( .A0(n25028), .A1(n24525), .B0(n25027), .Y(n2435) );
  OAI21XL U25804 ( .A0(n25030), .A1(n3057), .B0(n25029), .Y(n25031) );
  OAI21XL U25805 ( .A0(n25059), .A1(n25929), .B0(n25032), .Y(n25033) );
  AOI222XL U25806 ( .A0(n25623), .A1(n4710), .B0(n25822), .B1(w2[33]), .C0(
        w2[65]), .C1(in_valid_w2), .Y(n2169) );
  OAI21XL U25807 ( .A0(n25059), .A1(n25918), .B0(n25034), .Y(n25035) );
  AOI222XL U25808 ( .A0(n25596), .A1(n4710), .B0(n25822), .B1(w2[35]), .C0(
        w2[67]), .C1(in_valid_w2), .Y(n2171) );
  OAI21XL U25809 ( .A0(n25059), .A1(n26271), .B0(n25036), .Y(n25037) );
  AOI222XL U25810 ( .A0(n25566), .A1(n4710), .B0(n25822), .B1(w2[37]), .C0(
        w2[69]), .C1(in_valid_w2), .Y(n2173) );
  OAI21XL U25811 ( .A0(n25059), .A1(n25919), .B0(n25038), .Y(n25039) );
  AOI222XL U25812 ( .A0(n25545), .A1(n4710), .B0(n25822), .B1(w2[39]), .C0(
        w2[71]), .C1(in_valid_w2), .Y(n2175) );
  OAI21XL U25813 ( .A0(n25059), .A1(n26272), .B0(n25040), .Y(n25041) );
  AOI222XL U25814 ( .A0(n25518), .A1(n25292), .B0(n25822), .B1(w2[41]), .C0(
        w2[73]), .C1(in_valid_w2), .Y(n2177) );
  OAI21XL U25815 ( .A0(n25059), .A1(n26007), .B0(n25042), .Y(n25043) );
  AOI222XL U25816 ( .A0(n25495), .A1(n25292), .B0(n25822), .B1(w2[43]), .C0(
        w2[75]), .C1(in_valid_w2), .Y(n2179) );
  OAI21XL U25817 ( .A0(n25059), .A1(n26273), .B0(n25044), .Y(n25045) );
  AOI222XL U25818 ( .A0(n25472), .A1(n25292), .B0(n25822), .B1(w2[45]), .C0(
        w2[77]), .C1(in_valid_w2), .Y(n2181) );
  OAI21XL U25819 ( .A0(n25059), .A1(n25920), .B0(n25046), .Y(n25047) );
  AOI222XL U25820 ( .A0(n25448), .A1(n25292), .B0(n25822), .B1(w2[47]), .C0(
        w2[79]), .C1(in_valid_w2), .Y(n2183) );
  AOI222XL U25821 ( .A0(n25421), .A1(n4710), .B0(n25822), .B1(w2[49]), .C0(
        w2[81]), .C1(in_valid_w2), .Y(n2185) );
  OAI21XL U25822 ( .A0(n25059), .A1(n25922), .B0(n25048), .Y(n25049) );
  AOI222XL U25823 ( .A0(n25392), .A1(n25292), .B0(n25822), .B1(w2[51]), .C0(
        w2[83]), .C1(in_valid_w2), .Y(n2187) );
  OAI21XL U25824 ( .A0(n25059), .A1(n25924), .B0(n25050), .Y(n25051) );
  AOI222XL U25825 ( .A0(n25371), .A1(n25292), .B0(n25822), .B1(w2[53]), .C0(
        w2[85]), .C1(in_valid_w2), .Y(n2189) );
  OAI21XL U25826 ( .A0(n25059), .A1(n25923), .B0(n25052), .Y(n25053) );
  AOI222XL U25827 ( .A0(n25384), .A1(n25292), .B0(n25822), .B1(w2[52]), .C0(
        w2[84]), .C1(in_valid_w2), .Y(n2188) );
  OAI21XL U25828 ( .A0(n25059), .A1(n26035), .B0(n25054), .Y(n25055) );
  AOI222XL U25829 ( .A0(n25407), .A1(n4710), .B0(n25822), .B1(w2[50]), .C0(
        w2[82]), .C1(in_valid_w2), .Y(n2186) );
  AOI222XL U25830 ( .A0(n25435), .A1(n25292), .B0(n25822), .B1(w2[48]), .C0(
        w2[80]), .C1(in_valid_w2), .Y(n2184) );
  AOI222XL U25831 ( .A0(n25459), .A1(n4710), .B0(n25822), .B1(w2[46]), .C0(
        w2[78]), .C1(in_valid_w2), .Y(n2182) );
  OAI21XL U25832 ( .A0(n25059), .A1(n26034), .B0(n25056), .Y(n25057) );
  AOI222XL U25833 ( .A0(n25485), .A1(n25292), .B0(n25822), .B1(w2[44]), .C0(
        w2[76]), .C1(in_valid_w2), .Y(n2180) );
  OAI21XL U25834 ( .A0(n25059), .A1(n26033), .B0(n25058), .Y(n25060) );
  AOI222XL U25835 ( .A0(n25508), .A1(n25292), .B0(n25822), .B1(w2[42]), .C0(
        w2[74]), .C1(in_valid_w2), .Y(n2178) );
  OAI21XL U25836 ( .A0(n25059), .A1(n26283), .B0(n25061), .Y(n25062) );
  AOI222XL U25837 ( .A0(n25533), .A1(n25292), .B0(n25822), .B1(w2[40]), .C0(
        w2[72]), .C1(in_valid_w2), .Y(n2176) );
  OAI21XL U25838 ( .A0(n25059), .A1(n26040), .B0(n25063), .Y(n25064) );
  AOI222XL U25839 ( .A0(n25558), .A1(n4710), .B0(n25822), .B1(w2[38]), .C0(
        w2[70]), .C1(in_valid_w2), .Y(n2174) );
  OAI21XL U25840 ( .A0(n25059), .A1(n26281), .B0(n25065), .Y(n25066) );
  AOI222XL U25841 ( .A0(n25577), .A1(n25292), .B0(n25822), .B1(w2[36]), .C0(
        w2[68]), .C1(in_valid_w2), .Y(n2172) );
  OAI21XL U25842 ( .A0(n25059), .A1(n25930), .B0(n25067), .Y(n25068) );
  AOI222XL U25843 ( .A0(n25609), .A1(n25292), .B0(n25822), .B1(w2[34]), .C0(
        w2[66]), .C1(in_valid_w2), .Y(n2170) );
  AOI222XL U25844 ( .A0(n25677), .A1(n4710), .B0(in_valid_w2), .B1(w2[64]), 
        .C0(w2[32]), .C1(n25822), .Y(n2168) );
  INVXL U25845 ( .A(n25070), .Y(n25069) );
  OAI21XL U25846 ( .A0(n25832), .A1(n25069), .B0(n25829), .Y(n25073) );
  NOR3XL U25847 ( .A(n25832), .B(n25072), .C(n25070), .Y(n25071) );
  AOI21XL U25848 ( .A0(n25076), .A1(n3065), .B0(n25075), .Y(n25077) );
  OAI21XL U25849 ( .A0(w1[315]), .A1(n3226), .B0(n25079), .Y(n1988) );
  AOI222XL U25850 ( .A0(n25080), .A1(n3216), .B0(w1[315]), .B1(n4578), .C0(
        n3061), .C1(w1[347]), .Y(n2116) );
  OAI21XL U25851 ( .A0(n3117), .A1(n26413), .B0(n25081), .Y(n25082) );
  AOI21XL U25852 ( .A0(n25083), .A1(n3216), .B0(n25082), .Y(n2118) );
  AOI222XL U25853 ( .A0(n25090), .A1(n3216), .B0(w1[347]), .B1(n4578), .C0(
        n23088), .C1(w1[379]), .Y(n2117) );
  AOI21XL U25854 ( .A0(n25541), .A1(w1[379]), .B0(n25085), .Y(n1990) );
  OAI21XL U25855 ( .A0(w1[347]), .A1(n4572), .B0(n25086), .Y(n1989) );
  OAI21XL U25856 ( .A0(w1[155]), .A1(n3226), .B0(n25087), .Y(n1863) );
  AOI22XL U25857 ( .A0(n3028), .A1(w1[27]), .B0(w1[155]), .B1(in_valid_w1), 
        .Y(n25088) );
  OAI21XL U25858 ( .A0(n3117), .A1(n26332), .B0(n25088), .Y(n25089) );
  AOI21XL U25859 ( .A0(n21112), .A1(w1[251]), .B0(n25089), .Y(n1862) );
  AOI22XL U25860 ( .A0(n25090), .A1(n25664), .B0(y11[27]), .B1(n24958), .Y(
        n25091) );
  AOI21XL U25861 ( .A0(n25675), .A1(n25170), .B0(n25092), .Y(n2483) );
  INVXL U25862 ( .A(n25093), .Y(n25097) );
  OAI21XL U25863 ( .A0(n25095), .A1(n3057), .B0(n25094), .Y(n25096) );
  AOI21XL U25864 ( .A0(n25675), .A1(n25097), .B0(n25096), .Y(n2447) );
  AOI21XL U25865 ( .A0(n25220), .A1(n25100), .B0(n25219), .Y(n25101) );
  OAI2BB1X1 U25866 ( .A0N(n25107), .A1N(n23643), .B0(n25101), .Y(mul5_out[27])
         );
  INVXL U25867 ( .A(n25842), .Y(n25105) );
  OAI21XL U25868 ( .A0(n25103), .A1(n3057), .B0(n25102), .Y(n25104) );
  AOI21XL U25869 ( .A0(n25675), .A1(n25105), .B0(n25104), .Y(n2451) );
  OAI21XL U25870 ( .A0(n25671), .A1(n4571), .B0(n25110), .Y(n2125) );
  AOI222XL U25871 ( .A0(n25683), .A1(n3216), .B0(w1[317]), .B1(n4577), .C0(
        n23088), .C1(w1[349]), .Y(n2124) );
  AOI21XL U25872 ( .A0(n25113), .A1(n3216), .B0(n25112), .Y(n2126) );
  OAI21XL U25873 ( .A0(w1[349]), .A1(n4574), .B0(n25114), .Y(n1997) );
  AOI21XL U25874 ( .A0(n25541), .A1(w1[381]), .B0(n25116), .Y(n1998) );
  OAI21XL U25875 ( .A0(w1[157]), .A1(n4573), .B0(n25117), .Y(n1871) );
  OAI21XL U25876 ( .A0(n3117), .A1(n26333), .B0(n25118), .Y(n25119) );
  AOI21XL U25877 ( .A0(n25541), .A1(w1[253]), .B0(n25119), .Y(n1870) );
  AOI21XL U25878 ( .A0(n25224), .A1(n3216), .B0(n25122), .Y(n2106) );
  ADDHXL U25879 ( .A(n25124), .B(n25123), .CO(n25125), .S(n20797) );
  AOI21XL U25880 ( .A0(n25220), .A1(n25134), .B0(n25219), .Y(n25135) );
  OAI2BB1X1 U25881 ( .A0N(n25136), .A1N(n23643), .B0(n25135), .Y(mul5_out[30])
         );
  INVXL U25882 ( .A(n25138), .Y(n25137) );
  AOI22XL U25883 ( .A0(n3029), .A1(n25138), .B0(n25290), .B1(n25137), .Y(
        n25642) );
  INVXL U25884 ( .A(n25642), .Y(n25647) );
  AOI222XL U25885 ( .A0(n25647), .A1(n25292), .B0(in_valid_w2), .B1(weight2[0]), .C0(w2[64]), .C1(n25822), .Y(n2200) );
  AOI21XL U25886 ( .A0(data[97]), .A1(n4582), .B0(n25139), .Y(n1711) );
  AOI21XL U25887 ( .A0(data[98]), .A1(n4584), .B0(n25140), .Y(n1712) );
  AOI21XL U25888 ( .A0(data[99]), .A1(n4584), .B0(n25141), .Y(n1713) );
  AOI21XL U25889 ( .A0(data[100]), .A1(n4586), .B0(n25142), .Y(n1714) );
  AOI21XL U25890 ( .A0(data[101]), .A1(n4586), .B0(n25143), .Y(n1715) );
  AOI21XL U25891 ( .A0(data[102]), .A1(n4583), .B0(n25144), .Y(n1716) );
  AOI21XL U25892 ( .A0(data[103]), .A1(n4581), .B0(n25145), .Y(n1717) );
  AOI21XL U25893 ( .A0(data[104]), .A1(n4583), .B0(n25146), .Y(n1718) );
  AOI21XL U25894 ( .A0(data[105]), .A1(n4581), .B0(n25147), .Y(n1719) );
  AOI21XL U25895 ( .A0(data[106]), .A1(n4586), .B0(n25148), .Y(n1720) );
  AOI21XL U25896 ( .A0(data[107]), .A1(n4586), .B0(n25149), .Y(n1721) );
  AOI21XL U25897 ( .A0(data[108]), .A1(n4584), .B0(n25150), .Y(n1722) );
  AOI21XL U25898 ( .A0(data[109]), .A1(n4584), .B0(n25151), .Y(n1723) );
  AOI21XL U25899 ( .A0(data[110]), .A1(n4582), .B0(n25152), .Y(n1724) );
  AOI21XL U25900 ( .A0(data[111]), .A1(n4585), .B0(n25153), .Y(n1725) );
  AOI21XL U25901 ( .A0(data[112]), .A1(n4586), .B0(n25154), .Y(n1726) );
  AOI21XL U25902 ( .A0(data[113]), .A1(n4581), .B0(n25155), .Y(n1727) );
  AOI21XL U25903 ( .A0(data[114]), .A1(n4586), .B0(n4771), .Y(n1728) );
  AOI21XL U25904 ( .A0(data[116]), .A1(n4581), .B0(n25157), .Y(n1730) );
  AOI21XL U25905 ( .A0(data[117]), .A1(n4582), .B0(n25158), .Y(n1731) );
  AOI21XL U25906 ( .A0(n25220), .A1(n25160), .B0(n25219), .Y(n25161) );
  OAI2BB1X1 U25907 ( .A0N(n25162), .A1N(n23643), .B0(n25161), .Y(mul5_out[28])
         );
  OAI21XL U25908 ( .A0(n26302), .A1(n3045), .B0(n25164), .Y(n25165) );
  AOI21XL U25909 ( .A0(n25166), .A1(n25767), .B0(n25165), .Y(n2292) );
  OAI21XL U25910 ( .A0(mul5_out[27]), .A1(n5434), .B0(n25171), .Y(n2350) );
  OAI21XL U25911 ( .A0(n26410), .A1(n3045), .B0(n25172), .Y(n25173) );
  AOI21XL U25912 ( .A0(n25767), .A1(n25174), .B0(n25173), .Y(n2291) );
  AOI21XL U25913 ( .A0(n25754), .A1(n25678), .B0(n25177), .Y(n2349) );
  AOI21XL U25914 ( .A0(n25220), .A1(n25179), .B0(n25219), .Y(n25180) );
  OAI2BB1X1 U25915 ( .A0N(n25181), .A1N(n23643), .B0(n25180), .Y(mul5_out[26])
         );
  ADDHXL U25916 ( .A(n25184), .B(n25183), .CO(n24284), .S(n25185) );
  OAI21XL U25917 ( .A0(n26297), .A1(n3045), .B0(n25186), .Y(n25187) );
  AOI21XL U25918 ( .A0(n25679), .A1(n25796), .B0(n25187), .Y(n2290) );
  AOI21XL U25919 ( .A0(n25754), .A1(n25191), .B0(n25190), .Y(n2347) );
  OAI21XL U25920 ( .A0(n26411), .A1(n3045), .B0(n25193), .Y(n25194) );
  AOI21XL U25921 ( .A0(n25195), .A1(n25767), .B0(n25194), .Y(n2289) );
  AOI21XL U25922 ( .A0(n25754), .A1(n25199), .B0(n25198), .Y(n2345) );
  OAI21XL U25923 ( .A0(n26282), .A1(n3045), .B0(n25202), .Y(n25203) );
  AOI21XL U25924 ( .A0(n25204), .A1(n25796), .B0(n25203), .Y(n2288) );
  AOI21XL U25925 ( .A0(data[125]), .A1(n4585), .B0(n25211), .Y(n1739) );
  AOI21XL U25926 ( .A0(data[124]), .A1(n4583), .B0(n25212), .Y(n1738) );
  AOI21XL U25927 ( .A0(data[123]), .A1(n4582), .B0(n25214), .Y(n1737) );
  AOI21XL U25928 ( .A0(data[122]), .A1(n4586), .B0(n25215), .Y(n1736) );
  AOI21XL U25929 ( .A0(data[121]), .A1(n4585), .B0(n25217), .Y(n1735) );
  AOI21XL U25930 ( .A0(data[120]), .A1(n4583), .B0(n25218), .Y(n1734) );
  AOI222XL U25931 ( .A0(n25227), .A1(n25292), .B0(w2[56]), .B1(n25822), .C0(
        w2[88]), .C1(in_valid_w2), .Y(n2192) );
  OAI21XL U25932 ( .A0(w1[344]), .A1(n4573), .B0(n25225), .Y(n1977) );
  OAI21XL U25933 ( .A0(n25227), .A1(n25584), .B0(n25226), .Y(n2105) );
  AOI222XL U25934 ( .A0(n25712), .A1(n3216), .B0(w1[312]), .B1(n4578), .C0(
        n3061), .C1(w1[344]), .Y(n2104) );
  OAI21XL U25935 ( .A0(w1[313]), .A1(n3226), .B0(n25228), .Y(n1980) );
  NAND2XL U25936 ( .A(n25233), .B(data[31]), .Y(n25235) );
  MXI2XL U25937 ( .A(w2[95]), .B(w2[63]), .S0(n23973), .Y(n25242) );
  OAI21XL U25938 ( .A0(n3121), .A1(n25660), .B0(n25249), .Y(n2555) );
  OAI21XL U25939 ( .A0(n25665), .A1(n3226), .B0(n25250), .Y(n2133) );
  OAI21XL U25940 ( .A0(n25697), .A1(n3226), .B0(n25251), .Y(n2132) );
  AOI21XL U25941 ( .A0(n25659), .A1(n3216), .B0(n25253), .Y(n2134) );
  OAI21XL U25942 ( .A0(w1[351]), .A1(n4573), .B0(n25254), .Y(n2005) );
  AOI21XL U25943 ( .A0(temp2[31]), .A1(n2983), .B0(n25259), .Y(n25260) );
  OAI21XL U25944 ( .A0(n4582), .A1(n25660), .B0(n25260), .Y(n2618) );
  INVXL U25945 ( .A(n25722), .Y(n25264) );
  OAI21XL U25946 ( .A0(n25262), .A1(n3057), .B0(n25261), .Y(n25263) );
  AOI21XL U25947 ( .A0(n25675), .A1(n25264), .B0(n25263), .Y(n2445) );
  OAI21XL U25948 ( .A0(n25275), .A1(n6219), .B0(n3077), .Y(n25276) );
  NOR2XL U25949 ( .A(n25282), .B(n25281), .Y(n25283) );
  NAND2XL U25950 ( .A(n25286), .B(n25285), .Y(n25288) );
  AOI22XL U25951 ( .A0(n24617), .A1(n25291), .B0(n25290), .B1(n25289), .Y(
        n25337) );
  INVXL U25952 ( .A(n25337), .Y(n25367) );
  AOI222XL U25953 ( .A0(n25367), .A1(n4710), .B0(n25822), .B1(w2[86]), .C0(
        weight2[22]), .C1(in_valid_w2), .Y(n2222) );
  INVXL U25954 ( .A(n25293), .Y(mul5_out[1]) );
  OAI21XL U25955 ( .A0(n3045), .A1(n25898), .B0(n25295), .Y(n25296) );
  AOI211XL U25956 ( .A0(n25329), .A1(n25298), .B0(n25297), .C0(n25296), .Y(
        n2265) );
  OAI21XL U25957 ( .A0(n25742), .A1(n25711), .B0(n25302), .Y(n2136) );
  OAI21XL U25958 ( .A0(n25624), .A1(n3118), .B0(n25303), .Y(n2137) );
  OAI21XL U25959 ( .A0(n25610), .A1(n3118), .B0(n25304), .Y(n2138) );
  OAI21XL U25960 ( .A0(n25597), .A1(n3118), .B0(n25305), .Y(n2139) );
  OAI21XL U25961 ( .A0(n25578), .A1(n3118), .B0(n25306), .Y(n2140) );
  OAI21XL U25962 ( .A0(n25568), .A1(n3118), .B0(n25307), .Y(n2141) );
  OAI21XL U25963 ( .A0(n25739), .A1(n3118), .B0(n25309), .Y(n2142) );
  OAI21XL U25964 ( .A0(n25546), .A1(n3118), .B0(n25310), .Y(n2143) );
  OAI21XL U25965 ( .A0(n25520), .A1(n3118), .B0(n25312), .Y(n2145) );
  OAI21XL U25966 ( .A0(n25509), .A1(n3118), .B0(n25313), .Y(n2146) );
  OAI21XL U25967 ( .A0(n25496), .A1(n3118), .B0(n25314), .Y(n2147) );
  OAI21XL U25968 ( .A0(n25486), .A1(n3118), .B0(n25315), .Y(n2148) );
  OAI21XL U25969 ( .A0(n25736), .A1(n3118), .B0(n25317), .Y(n2149) );
  OAI21XL U25970 ( .A0(n25460), .A1(n3118), .B0(n25318), .Y(n2150) );
  OAI21XL U25971 ( .A0(n25734), .A1(n25711), .B0(n25320), .Y(n2151) );
  OAI21XL U25972 ( .A0(n25436), .A1(n25711), .B0(n25321), .Y(n2152) );
  OAI21XL U25973 ( .A0(n25422), .A1(n25711), .B0(n25322), .Y(n2153) );
  OAI21XL U25974 ( .A0(n25732), .A1(n25711), .B0(n25324), .Y(n2154) );
  OAI21XL U25975 ( .A0(n25393), .A1(n25711), .B0(n25325), .Y(n2155) );
  OAI21XL U25976 ( .A0(n25385), .A1(n25711), .B0(n25326), .Y(n2156) );
  OAI21XL U25977 ( .A0(n25372), .A1(n25711), .B0(n25327), .Y(n2157) );
  OAI21XL U25978 ( .A0(n3045), .A1(n25909), .B0(n25332), .Y(n25333) );
  AOI211XL U25979 ( .A0(n25335), .A1(n4950), .B0(n25334), .C0(n25333), .Y(
        n2264) );
  INVXL U25980 ( .A(n25747), .Y(n25339) );
  AOI22XL U25981 ( .A0(n25025), .A1(y12[22]), .B0(n3122), .B1(y11[22]), .Y(
        n25336) );
  OAI21XL U25982 ( .A0(n25337), .A1(n3057), .B0(n25336), .Y(n25338) );
  NOR2XL U25983 ( .A(n25340), .B(n3075), .Y(n25351) );
  NAND2XL U25984 ( .A(n3030), .B(n25344), .Y(n25345) );
  OAI21XL U25985 ( .A0(n25347), .A1(n6177), .B0(n3075), .Y(n25348) );
  NOR2XL U25986 ( .A(n25354), .B(n25353), .Y(n25355) );
  NAND2XL U25987 ( .A(n25358), .B(n25357), .Y(n25360) );
  XOR2X1 U25988 ( .A(n25360), .B(n25359), .Y(n25361) );
  AOI222XL U25989 ( .A0(n25824), .A1(n3216), .B0(w1[310]), .B1(n4576), .C0(
        n3061), .C1(w1[342]), .Y(n2096) );
  AOI21XL U25990 ( .A0(n25367), .A1(n3216), .B0(n25366), .Y(n2098) );
  OAI21XL U25991 ( .A0(w1[342]), .A1(n25584), .B0(n25368), .Y(n1969) );
  OAI21XL U25992 ( .A0(w1[214]), .A1(n25584), .B0(n25369), .Y(n1841) );
  AOI222XL U25993 ( .A0(n25372), .A1(n3216), .B0(w1[309]), .B1(n4576), .C0(
        n23088), .C1(w1[341]), .Y(n2092) );
  INVXL U25994 ( .A(n25373), .Y(n25376) );
  AOI21XL U25995 ( .A0(n25376), .A1(n3216), .B0(n25375), .Y(n2094) );
  OAI21XL U25996 ( .A0(w1[341]), .A1(n25584), .B0(n25377), .Y(n1965) );
  AOI22XL U25997 ( .A0(n25378), .A1(n25638), .B0(n2983), .B1(temp2[20]), .Y(
        n25381) );
  NAND2XL U25998 ( .A(n25379), .B(n25636), .Y(n25380) );
  OAI211XL U25999 ( .A0(n25382), .A1(n4581), .B0(n25381), .C0(n25380), .Y(
        n2577) );
  AOI222XL U26000 ( .A0(n25385), .A1(n3216), .B0(w1[308]), .B1(n4576), .C0(
        n23088), .C1(w1[340]), .Y(n2088) );
  INVXL U26001 ( .A(n25386), .Y(n25389) );
  AOI21XL U26002 ( .A0(n25389), .A1(n3216), .B0(n25388), .Y(n2090) );
  OAI21XL U26003 ( .A0(w1[340]), .A1(n25584), .B0(n25390), .Y(n1961) );
  AOI222XL U26004 ( .A0(n25393), .A1(n3216), .B0(w1[307]), .B1(n4576), .C0(
        n3061), .C1(w1[339]), .Y(n2084) );
  INVXL U26005 ( .A(n25394), .Y(n25397) );
  AOI21XL U26006 ( .A0(n25397), .A1(n3216), .B0(n25396), .Y(n2086) );
  OAI21XL U26007 ( .A0(w1[339]), .A1(n3226), .B0(n25398), .Y(n1957) );
  OAI21XL U26008 ( .A0(w1[275]), .A1(n25584), .B0(n25399), .Y(n1959) );
  AOI21XL U26009 ( .A0(n25541), .A1(w1[371]), .B0(n25401), .Y(n1958) );
  OAI21XL U26010 ( .A0(w1[211]), .A1(n4571), .B0(n25402), .Y(n1829) );
  OAI21XL U26011 ( .A0(w1[179]), .A1(n3226), .B0(n25403), .Y(n1828) );
  AOI21XL U26012 ( .A0(n25541), .A1(w1[243]), .B0(n25405), .Y(n1830) );
  AOI222XL U26013 ( .A0(n25732), .A1(n3216), .B0(w1[306]), .B1(n25410), .C0(
        n23088), .C1(w1[338]), .Y(n2080) );
  INVXL U26014 ( .A(n25408), .Y(n25412) );
  AOI21XL U26015 ( .A0(n25412), .A1(n3216), .B0(n25411), .Y(n2082) );
  OAI21XL U26016 ( .A0(w1[338]), .A1(n4571), .B0(n25413), .Y(n1953) );
  OAI21XL U26017 ( .A0(w1[306]), .A1(n4572), .B0(n25414), .Y(n1952) );
  AOI21XL U26018 ( .A0(n21112), .A1(w1[370]), .B0(n25416), .Y(n1954) );
  OAI21XL U26019 ( .A0(w1[210]), .A1(n4571), .B0(n25417), .Y(n1825) );
  AOI21XL U26020 ( .A0(n25541), .A1(w1[242]), .B0(n25419), .Y(n1826) );
  AOI222XL U26021 ( .A0(n25422), .A1(n3216), .B0(w1[305]), .B1(n4578), .C0(
        n23088), .C1(w1[337]), .Y(n2076) );
  INVXL U26022 ( .A(n25423), .Y(n25426) );
  AOI21XL U26023 ( .A0(n25426), .A1(n3216), .B0(n25425), .Y(n2078) );
  OAI21XL U26024 ( .A0(w1[337]), .A1(n4572), .B0(n25427), .Y(n1949) );
  AOI21XL U26025 ( .A0(n25541), .A1(w1[369]), .B0(n25430), .Y(n1950) );
  OAI21XL U26026 ( .A0(w1[145]), .A1(n4572), .B0(n25431), .Y(n1823) );
  OAI21XL U26027 ( .A0(n3117), .A1(n26338), .B0(n25432), .Y(n25433) );
  AOI21XL U26028 ( .A0(n25541), .A1(w1[241]), .B0(n25433), .Y(n1822) );
  AOI222XL U26029 ( .A0(n25436), .A1(n3216), .B0(w1[304]), .B1(n4577), .C0(
        n3061), .C1(w1[336]), .Y(n2072) );
  INVXL U26030 ( .A(n25437), .Y(n25440) );
  AOI21XL U26031 ( .A0(n25440), .A1(n3216), .B0(n25439), .Y(n2074) );
  OAI21XL U26032 ( .A0(w1[272]), .A1(n4571), .B0(n25441), .Y(n1947) );
  OAI21XL U26033 ( .A0(n3117), .A1(n26327), .B0(n25442), .Y(n25443) );
  AOI21XL U26034 ( .A0(n25541), .A1(w1[368]), .B0(n25443), .Y(n1946) );
  OAI21XL U26035 ( .A0(w1[176]), .A1(n4572), .B0(n25444), .Y(n1816) );
  OAI21XL U26036 ( .A0(n3117), .A1(n26339), .B0(n25445), .Y(n25446) );
  AOI21XL U26037 ( .A0(n25541), .A1(w1[240]), .B0(n25446), .Y(n1818) );
  AOI222XL U26038 ( .A0(n25734), .A1(n3216), .B0(w1[303]), .B1(n4577), .C0(
        n3061), .C1(w1[335]), .Y(n2068) );
  INVXL U26039 ( .A(n25449), .Y(n25452) );
  AOI21XL U26040 ( .A0(n25452), .A1(n3216), .B0(n25451), .Y(n2070) );
  OAI21XL U26041 ( .A0(w1[335]), .A1(n4572), .B0(n25453), .Y(n1941) );
  AOI21XL U26042 ( .A0(n25541), .A1(w1[367]), .B0(n25455), .Y(n1942) );
  OAI21XL U26043 ( .A0(n3117), .A1(n26340), .B0(n25456), .Y(n25457) );
  AOI21XL U26044 ( .A0(n25541), .A1(w1[239]), .B0(n25457), .Y(n1814) );
  AOI222XL U26045 ( .A0(n25460), .A1(n3216), .B0(w1[302]), .B1(n4576), .C0(
        n3061), .C1(w1[334]), .Y(n2064) );
  INVXL U26046 ( .A(n25461), .Y(n25464) );
  AOI21XL U26047 ( .A0(n25464), .A1(n3216), .B0(n25463), .Y(n2066) );
  OAI21XL U26048 ( .A0(w1[334]), .A1(n4573), .B0(n25465), .Y(n1937) );
  AOI21XL U26049 ( .A0(n21112), .A1(w1[366]), .B0(n25467), .Y(n1938) );
  OAI21XL U26050 ( .A0(w1[142]), .A1(n4572), .B0(n25468), .Y(n1811) );
  OAI21XL U26051 ( .A0(n3117), .A1(n26341), .B0(n25469), .Y(n25470) );
  AOI21XL U26052 ( .A0(n25541), .A1(w1[238]), .B0(n25470), .Y(n1810) );
  AOI222XL U26053 ( .A0(n25736), .A1(n3216), .B0(w1[301]), .B1(n4576), .C0(
        n3061), .C1(w1[333]), .Y(n2060) );
  INVXL U26054 ( .A(n25473), .Y(n25476) );
  AOI21XL U26055 ( .A0(n25476), .A1(n21112), .B0(n25475), .Y(n2062) );
  OAI21XL U26056 ( .A0(w1[333]), .A1(n4573), .B0(n25477), .Y(n1933) );
  OAI21XL U26057 ( .A0(w1[301]), .A1(n4573), .B0(n25478), .Y(n1932) );
  AOI21XL U26058 ( .A0(n21112), .A1(w1[365]), .B0(n25480), .Y(n1934) );
  OAI21XL U26059 ( .A0(n3117), .A1(n26342), .B0(n25481), .Y(n25482) );
  AOI21XL U26060 ( .A0(n25541), .A1(w1[237]), .B0(n25482), .Y(n1806) );
  OAI222XL U26061 ( .A0(n3226), .A1(n25486), .B0(n3228), .B1(w1[332]), .C0(
        n3117), .C1(w1[300]), .Y(n2056) );
  INVXL U26062 ( .A(n25487), .Y(n25490) );
  AOI21XL U26063 ( .A0(n25490), .A1(n3216), .B0(n25489), .Y(n2058) );
  OAI21XL U26064 ( .A0(w1[332]), .A1(n4571), .B0(n25491), .Y(n1929) );
  OAI21XL U26065 ( .A0(w1[172]), .A1(n4573), .B0(n25492), .Y(n1800) );
  OAI21XL U26066 ( .A0(w1[140]), .A1(n4573), .B0(n25493), .Y(n1803) );
  AOI222XL U26067 ( .A0(n25496), .A1(n3216), .B0(w1[299]), .B1(n4578), .C0(
        n23088), .C1(w1[331]), .Y(n2052) );
  INVXL U26068 ( .A(n25497), .Y(n25500) );
  AOI21XL U26069 ( .A0(n25500), .A1(n3216), .B0(n25499), .Y(n2054) );
  OAI21XL U26070 ( .A0(w1[331]), .A1(n4574), .B0(n25501), .Y(n1925) );
  AOI22XL U26071 ( .A0(n25502), .A1(n25636), .B0(n2983), .B1(temp2[10]), .Y(
        n25505) );
  NAND2XL U26072 ( .A(n25503), .B(n25638), .Y(n25504) );
  OAI211XL U26073 ( .A0(n25506), .A1(n4582), .B0(n25505), .C0(n25504), .Y(
        n2597) );
  AOI222XL U26074 ( .A0(n25509), .A1(n3216), .B0(w1[298]), .B1(n3052), .C0(
        n3061), .C1(w1[330]), .Y(n2048) );
  INVXL U26075 ( .A(n25510), .Y(n25513) );
  AOI21XL U26076 ( .A0(n25513), .A1(n3216), .B0(n25512), .Y(n2050) );
  OAI21XL U26077 ( .A0(w1[330]), .A1(n4573), .B0(n25514), .Y(n1921) );
  OAI21XL U26078 ( .A0(w1[266]), .A1(n4572), .B0(n25515), .Y(n1923) );
  OAI21XL U26079 ( .A0(w1[170]), .A1(n4574), .B0(n25516), .Y(n1792) );
  OAI21XL U26080 ( .A0(n25520), .A1(n3226), .B0(n25519), .Y(n2044) );
  INVXL U26081 ( .A(n25521), .Y(n25524) );
  AOI21XL U26082 ( .A0(n25524), .A1(n3216), .B0(n25523), .Y(n2046) );
  OAI21XL U26083 ( .A0(w1[329]), .A1(n4574), .B0(n25525), .Y(n1917) );
  OAI21XL U26084 ( .A0(w1[265]), .A1(n25584), .B0(n25526), .Y(n1919) );
  AOI22XL U26085 ( .A0(n25527), .A1(n25636), .B0(n2984), .B1(temp2[8]), .Y(
        n25530) );
  NAND2XL U26086 ( .A(n25528), .B(n25638), .Y(n25529) );
  OAI211XL U26087 ( .A0(n25531), .A1(n4582), .B0(n25530), .C0(n25529), .Y(
        n2601) );
  INVXL U26088 ( .A(n25536), .Y(n25539) );
  AOI21XL U26089 ( .A0(n25539), .A1(n3216), .B0(n25538), .Y(n2042) );
  OAI21XL U26090 ( .A0(w1[328]), .A1(n4574), .B0(n25540), .Y(n1913) );
  OAI21XL U26091 ( .A0(w1[264]), .A1(n4573), .B0(n25543), .Y(n1915) );
  AOI222XL U26092 ( .A0(n25546), .A1(n3216), .B0(w1[295]), .B1(n4576), .C0(
        n3061), .C1(w1[327]), .Y(n2036) );
  INVXL U26093 ( .A(n25547), .Y(n25550) );
  AOI21XL U26094 ( .A0(n25550), .A1(n3216), .B0(n25549), .Y(n2038) );
  OAI21XL U26095 ( .A0(w1[327]), .A1(n3226), .B0(n25551), .Y(n1909) );
  AOI22XL U26096 ( .A0(n25552), .A1(n25636), .B0(n2983), .B1(temp2[6]), .Y(
        n25555) );
  NAND2XL U26097 ( .A(n25553), .B(n25638), .Y(n25554) );
  OAI211XL U26098 ( .A0(n25556), .A1(n4586), .B0(n25555), .C0(n25554), .Y(
        n2605) );
  AOI222XL U26099 ( .A0(n25739), .A1(n3216), .B0(w1[294]), .B1(n4578), .C0(
        n3061), .C1(w1[326]), .Y(n2032) );
  INVXL U26100 ( .A(n25559), .Y(n25562) );
  AOI21XL U26101 ( .A0(n25562), .A1(n3216), .B0(n25561), .Y(n2034) );
  OAI21XL U26102 ( .A0(w1[326]), .A1(n3226), .B0(n25563), .Y(n1905) );
  OAI21XL U26103 ( .A0(w1[198]), .A1(n25584), .B0(n25564), .Y(n1777) );
  AOI222XL U26104 ( .A0(n25568), .A1(n3216), .B0(w1[293]), .B1(n4578), .C0(
        n23088), .C1(w1[325]), .Y(n2028) );
  INVXL U26105 ( .A(n25569), .Y(n25572) );
  AOI21XL U26106 ( .A0(n25572), .A1(n3216), .B0(n25571), .Y(n2030) );
  OAI21XL U26107 ( .A0(w1[325]), .A1(n25584), .B0(n25573), .Y(n1901) );
  OAI21XL U26108 ( .A0(w1[197]), .A1(n25584), .B0(n25574), .Y(n1773) );
  OAI21XL U26109 ( .A0(w1[133]), .A1(n3226), .B0(n25575), .Y(n1775) );
  AOI222XL U26110 ( .A0(n25578), .A1(n3216), .B0(w1[292]), .B1(n4578), .C0(
        n3061), .C1(w1[324]), .Y(n2024) );
  INVXL U26111 ( .A(n25579), .Y(n25582) );
  AOI21XL U26112 ( .A0(n25582), .A1(n3216), .B0(n25581), .Y(n2026) );
  OAI21XL U26113 ( .A0(w1[324]), .A1(n25584), .B0(n25583), .Y(n1897) );
  AOI21XL U26114 ( .A0(n25541), .A1(w1[356]), .B0(n25586), .Y(n1898) );
  OAI21XL U26115 ( .A0(w1[196]), .A1(n3226), .B0(n25587), .Y(n1769) );
  AOI21XL U26116 ( .A0(n25541), .A1(w1[228]), .B0(n25589), .Y(n1770) );
  AOI22XL U26117 ( .A0(n25590), .A1(n25636), .B0(n2984), .B1(temp2[3]), .Y(
        n25593) );
  NAND2XL U26118 ( .A(n25591), .B(n25638), .Y(n25592) );
  OAI211XL U26119 ( .A0(n25594), .A1(n4585), .B0(n25593), .C0(n25592), .Y(
        n2611) );
  AOI222XL U26120 ( .A0(n25597), .A1(n3216), .B0(w1[291]), .B1(n4577), .C0(
        n23088), .C1(w1[323]), .Y(n2020) );
  INVXL U26121 ( .A(n25598), .Y(n25601) );
  AOI21XL U26122 ( .A0(n25601), .A1(n3216), .B0(n25600), .Y(n2022) );
  OAI21XL U26123 ( .A0(w1[323]), .A1(n3226), .B0(n25602), .Y(n1893) );
  AOI21XL U26124 ( .A0(n25541), .A1(w1[355]), .B0(n25604), .Y(n1894) );
  OAI21XL U26125 ( .A0(w1[131]), .A1(n3226), .B0(n25605), .Y(n1767) );
  OAI21XL U26126 ( .A0(n3117), .A1(n26349), .B0(n25606), .Y(n25607) );
  AOI21XL U26127 ( .A0(n21112), .A1(w1[227]), .B0(n25607), .Y(n1766) );
  AOI222XL U26128 ( .A0(n25610), .A1(n3216), .B0(w1[290]), .B1(n4578), .C0(
        n3061), .C1(w1[322]), .Y(n2016) );
  INVXL U26129 ( .A(n25611), .Y(n25614) );
  AOI21XL U26130 ( .A0(n25614), .A1(n3216), .B0(n25613), .Y(n2018) );
  OAI21XL U26131 ( .A0(w1[322]), .A1(n3226), .B0(n25615), .Y(n1889) );
  OAI21XL U26132 ( .A0(w1[290]), .A1(n4574), .B0(n25616), .Y(n1888) );
  AOI21XL U26133 ( .A0(n25541), .A1(w1[354]), .B0(n25618), .Y(n1890) );
  OAI21XL U26134 ( .A0(w1[130]), .A1(n25584), .B0(n25619), .Y(n1763) );
  OAI21XL U26135 ( .A0(n3117), .A1(n26350), .B0(n25620), .Y(n25621) );
  AOI21XL U26136 ( .A0(n25541), .A1(w1[226]), .B0(n25621), .Y(n1762) );
  AOI222XL U26137 ( .A0(n25624), .A1(n3216), .B0(w1[289]), .B1(n4578), .C0(
        n23088), .C1(w1[321]), .Y(n2012) );
  INVXL U26138 ( .A(n25625), .Y(n25628) );
  AOI21XL U26139 ( .A0(n25628), .A1(n3216), .B0(n25627), .Y(n2014) );
  OAI21XL U26140 ( .A0(w1[321]), .A1(n4573), .B0(n25629), .Y(n1885) );
  AOI21XL U26141 ( .A0(n25541), .A1(w1[353]), .B0(n25631), .Y(n1886) );
  OAI21XL U26142 ( .A0(w1[193]), .A1(n4572), .B0(n25632), .Y(n1757) );
  AOI21XL U26143 ( .A0(n25541), .A1(w1[225]), .B0(n25634), .Y(n1758) );
  AOI22XL U26144 ( .A0(n25636), .A1(n25635), .B0(n2983), .B1(temp2[0]), .Y(
        n25640) );
  NAND2XL U26145 ( .A(n25638), .B(n25637), .Y(n25639) );
  AOI22XL U26146 ( .A0(n24739), .A1(y12[0]), .B0(n3122), .B1(y11[0]), .Y(
        n25641) );
  OAI21XL U26147 ( .A0(n25642), .A1(n3057), .B0(n25641), .Y(n25643) );
  AOI21XL U26148 ( .A0(n25644), .A1(n25675), .B0(n25643), .Y(n2393) );
  AOI21XL U26149 ( .A0(n25647), .A1(n3216), .B0(n25646), .Y(n2010) );
  AOI21XL U26150 ( .A0(n25541), .A1(w1[352]), .B0(n25649), .Y(n1882) );
  OAI21XL U26151 ( .A0(w1[320]), .A1(n4571), .B0(n25650), .Y(n1881) );
  OAI21XL U26152 ( .A0(w1[288]), .A1(n4571), .B0(n25651), .Y(n1880) );
  OAI21XL U26153 ( .A0(w1[192]), .A1(n4574), .B0(n25652), .Y(n1753) );
  OAI21XL U26154 ( .A0(w1[128]), .A1(n4574), .B0(n25653), .Y(n1755) );
  AOI21XL U26155 ( .A0(n25541), .A1(w1[224]), .B0(n25655), .Y(n1754) );
  OAI21XL U26156 ( .A0(n25660), .A1(n25693), .B0(n25657), .Y(n25658) );
  AOI21XL U26157 ( .A0(n25659), .A1(n3025), .B0(n25658), .Y(n2455) );
  OAI21XL U26158 ( .A0(n25693), .A1(n25670), .B0(n25662), .Y(n25663) );
  AOI21XL U26159 ( .A0(n25665), .A1(n25664), .B0(n25663), .Y(n2487) );
  OAI21XL U26160 ( .A0(n4584), .A1(n25670), .B0(n25669), .Y(n2619) );
  AOI22XL U26161 ( .A0(n25671), .A1(n3025), .B0(y11[29]), .B1(n24958), .Y(
        n25672) );
  AOI21XL U26162 ( .A0(n25675), .A1(n25674), .B0(n25673), .Y(n2485) );
  AOI222XL U26163 ( .A0(n25742), .A1(n3216), .B0(w1[288]), .B1(n4577), .C0(
        n23088), .C1(w1[320]), .Y(n2008) );
  INVXL U26164 ( .A(n25678), .Y(n25681) );
  OAI21XL U26165 ( .A0(n25697), .A1(n25711), .B0(n25682), .Y(n2167) );
  INVXL U26166 ( .A(n25683), .Y(n25685) );
  AOI22XL U26167 ( .A0(n24739), .A1(y10[29]), .B0(n3122), .B1(y12[29]), .Y(
        n25684) );
  AOI21XL U26168 ( .A0(n25840), .A1(n24525), .B0(n25686), .Y(n2450) );
  AOI22XL U26169 ( .A0(n25815), .A1(y10[0]), .B0(n3122), .B1(y12[0]), .Y(
        n25688) );
  OAI21XL U26170 ( .A0(n25689), .A1(n3057), .B0(n25688), .Y(n25690) );
  AOI21XL U26171 ( .A0(n25745), .A1(n6161), .B0(n25690), .Y(n2392) );
  AOI22XL U26172 ( .A0(n25025), .A1(y10[31]), .B0(n3122), .B1(y12[31]), .Y(
        n25692) );
  OAI21XL U26173 ( .A0(n25694), .A1(n25693), .B0(n25692), .Y(n25695) );
  AOI21XL U26174 ( .A0(n25697), .A1(n25696), .B0(n25695), .Y(n2454) );
  OAI21XL U26175 ( .A0(w1[350]), .A1(n4574), .B0(n25698), .Y(n2001) );
  AOI21XL U26176 ( .A0(n25704), .A1(n25703), .B0(n25702), .Y(n25705) );
  AOI21XL U26177 ( .A0(n25707), .A1(n3065), .B0(n25706), .Y(n25708) );
  OAI21XL U26178 ( .A0(n25832), .A1(n25713), .B0(n25829), .Y(n25717) );
  INVXL U26179 ( .A(n25713), .Y(n25714) );
  NOR3XL U26180 ( .A(n25832), .B(n25716), .C(n25714), .Y(n25715) );
  AOI21XL U26181 ( .A0(n25720), .A1(n3065), .B0(n25719), .Y(n25721) );
  AOI22XL U26182 ( .A0(n25725), .A1(n25724), .B0(n25723), .B1(temp0[21]), .Y(
        n25726) );
  AOI222XL U26183 ( .A0(n25733), .A1(n25737), .B0(n25743), .B1(y20[18]), .C0(
        n25732), .C1(n20890), .Y(n2378) );
  AOI222XL U26184 ( .A0(n25738), .A1(n25737), .B0(n25743), .B1(y20[13]), .C0(
        n25736), .C1(n20890), .Y(n2373) );
  AOI22XL U26185 ( .A0(n25821), .A1(n25664), .B0(y11[22]), .B1(n25815), .Y(
        n25746) );
  AOI21XL U26186 ( .A0(n3060), .A1(n25749), .B0(n25748), .Y(n2478) );
  AOI21XL U26187 ( .A0(n25754), .A1(n25753), .B0(n25752), .Y(n2339) );
  AOI211XL U26188 ( .A0(n25762), .A1(n25761), .B0(n25760), .C0(n25759), .Y(
        n2341) );
  OAI21XL U26189 ( .A0(n3045), .A1(n25915), .B0(n25765), .Y(n25766) );
  OAI21XL U26190 ( .A0(n26412), .A1(n3045), .B0(n25768), .Y(n25769) );
  AOI21XL U26191 ( .A0(n25813), .A1(n25770), .B0(n25769), .Y(n2293) );
  AOI21XL U26192 ( .A0(n25754), .A1(n25803), .B0(n25772), .Y(n2343) );
  NAND2XL U26193 ( .A(n24031), .B(n25775), .Y(n25781) );
  ADDHXL U26194 ( .A(n25773), .B(n25774), .CO(n25776), .S(n24032) );
  NAND2XL U26195 ( .A(n25778), .B(n25777), .Y(n25780) );
  AOI21XL U26196 ( .A0(n25754), .A1(n25819), .B0(n25784), .Y(n2357) );
  ADDHXL U26197 ( .A(n25788), .B(n25789), .CO(n25790), .S(n24051) );
  AOI21XL U26198 ( .A0(n24048), .A1(n25791), .B0(n3004), .Y(n25792) );
  OAI2BB1X1 U26199 ( .A0N(n3005), .A1N(n25793), .B0(n25792), .Y(n25797) );
  OAI21XL U26200 ( .A0(n26303), .A1(n3045), .B0(n25794), .Y(n25795) );
  AOI21XL U26201 ( .A0(n25796), .A1(n25797), .B0(n25795), .Y(n2294) );
  INVXL U26202 ( .A(n25819), .Y(n25799) );
  OAI21XL U26203 ( .A0(n25816), .A1(n4574), .B0(n25800), .Y(n2129) );
  AOI222XL U26204 ( .A0(n25801), .A1(n3216), .B0(w1[318]), .B1(n4577), .C0(
        n3061), .C1(w1[350]), .Y(n2128) );
  OAI21XL U26205 ( .A0(w1[318]), .A1(n4572), .B0(n25802), .Y(n2000) );
  INVXL U26206 ( .A(n25803), .Y(n25809) );
  AOI21XL U26207 ( .A0(n24048), .A1(n25804), .B0(n3004), .Y(n25805) );
  OAI2BB1X1 U26208 ( .A0N(n3005), .A1N(n25806), .B0(n25805), .Y(n25814) );
  AOI222XL U26209 ( .A0(n25810), .A1(n25292), .B0(w2[55]), .B1(n25822), .C0(
        w2[87]), .C1(in_valid_w2), .Y(n2191) );
  OAI21XL U26210 ( .A0(n26286), .A1(n3045), .B0(n25811), .Y(n25812) );
  AOI21XL U26211 ( .A0(n25813), .A1(n25814), .B0(n25812), .Y(n2287) );
  AOI22XL U26212 ( .A0(n25816), .A1(n25664), .B0(y11[30]), .B1(n25815), .Y(
        n25817) );
  AOI21XL U26213 ( .A0(n3060), .A1(n25819), .B0(n25818), .Y(n2486) );
  AOI222XL U26214 ( .A0(n25821), .A1(n4710), .B0(n25820), .B1(w2[54]), .C0(
        w2[86]), .C1(in_valid_w2), .Y(n2190) );
  OAI21XL U26215 ( .A0(n25824), .A1(n25711), .B0(n25823), .Y(n2158) );
  AOI22XL U26216 ( .A0(n25815), .A1(y10[22]), .B0(n3122), .B1(y12[22]), .Y(
        n25825) );
  OAI21XL U26217 ( .A0(n25826), .A1(n3057), .B0(n25825), .Y(n25827) );
  AOI21XL U26218 ( .A0(n25828), .A1(n6161), .B0(n25827), .Y(n2436) );
  INVXL U26219 ( .A(n25831), .Y(n25830) );
  OAI21XL U26220 ( .A0(n25832), .A1(n25830), .B0(n25829), .Y(n25836) );
  NOR3XL U26221 ( .A(n25832), .B(n25835), .C(n25831), .Y(n25833) );
  AOI21XL U26222 ( .A0(n25840), .A1(in_valid_d), .B0(n25839), .Y(n25841) );
  AOI21XL U26223 ( .A0(n25845), .A1(n25541), .B0(n25844), .Y(n2130) );
  AOI21XL U26224 ( .A0(n25541), .A1(w1[382]), .B0(n25847), .Y(n2002) );
  OAI21XL U26225 ( .A0(n3117), .A1(n26351), .B0(n25849), .Y(n25850) );
  AOI21XL U26226 ( .A0(n25541), .A1(w1[254]), .B0(n25850), .Y(n1874) );
  INVXL U26227 ( .A(n25851), .Y(n25855) );
  AOI22XL U26228 ( .A0(n24739), .A1(y12[30]), .B0(n3122), .B1(y11[30]), .Y(
        n25852) );
  OAI21XL U26229 ( .A0(n25853), .A1(n3057), .B0(n25852), .Y(n25854) );
  AOI21XL U26230 ( .A0(n3060), .A1(n25855), .B0(n25854), .Y(n2453) );
  AOI21XL U26231 ( .A0(iter[8]), .A1(n25858), .B0(n25856), .Y(n25857) );
  OAI21XL U26232 ( .A0(iter[8]), .A1(n25858), .B0(n25857), .Y(n1749) );
  CMPR42X1 U26233 ( .A(M6_mult_x_15_n1167), .B(M6_mult_x_15_n588), .C(
        M6_mult_x_15_n585), .D(M6_mult_x_15_n595), .ICI(M6_mult_x_15_n591), 
        .S(M6_mult_x_15_n582), .ICO(M6_mult_x_15_n580), .CO(M6_mult_x_15_n581)
         );
  CMPR42X1 U26234 ( .A(M6_mult_x_15_n1156), .B(M6_mult_x_15_n1180), .C(
        M6_mult_x_15_n707), .D(M6_mult_x_15_n1204), .ICI(M6_mult_x_15_n710), 
        .S(M6_mult_x_15_n705), .ICO(M6_mult_x_15_n703), .CO(M6_mult_x_15_n704)
         );
  CMPR42X1 U26235 ( .A(M6_mult_x_15_n1115), .B(M6_mult_x_15_n544), .C(
        M6_mult_x_15_n551), .D(M6_mult_x_15_n541), .ICI(M6_mult_x_15_n547), 
        .S(M6_mult_x_15_n538), .ICO(M6_mult_x_15_n536), .CO(M6_mult_x_15_n537)
         );
  CMPR42X1 U26236 ( .A(M6_mult_x_15_n1194), .B(M6_mult_x_15_n627), .C(
        M6_mult_x_15_n628), .D(M6_mult_x_15_n618), .ICI(M6_mult_x_15_n624), 
        .S(M6_mult_x_15_n615), .ICO(M6_mult_x_15_n613), .CO(M6_mult_x_15_n614)
         );
  CMPR42X1 U26237 ( .A(M6_mult_x_15_n1137), .B(M6_mult_x_15_n1065), .C(
        M6_mult_x_15_n1089), .D(M6_mult_x_15_n1113), .ICI(M6_mult_x_15_n524), 
        .S(M6_mult_x_15_n521), .ICO(M6_mult_x_15_n519), .CO(M6_mult_x_15_n520)
         );
  CMPR42X1 U26238 ( .A(M6_mult_x_15_n1070), .B(M6_mult_x_15_n1094), .C(
        M6_mult_x_15_n1166), .D(M6_mult_x_15_n586), .ICI(M6_mult_x_15_n1142), 
        .S(M6_mult_x_15_n574), .ICO(M6_mult_x_15_n572), .CO(M6_mult_x_15_n573)
         );
  CMPR42X1 U26239 ( .A(M6_mult_x_15_n1122), .B(M6_mult_x_15_n1146), .C(
        M6_mult_x_15_n1170), .D(M6_mult_x_15_n631), .ICI(M6_mult_x_15_n621), 
        .S(M6_mult_x_15_n618), .ICO(M6_mult_x_15_n616), .CO(M6_mult_x_15_n617)
         );
  CMPR42X1 U26240 ( .A(M6_mult_x_15_n1145), .B(M6_mult_x_15_n1121), .C(
        M6_mult_x_15_n1193), .D(M6_mult_x_15_n1169), .ICI(M6_mult_x_15_n616), 
        .S(M6_mult_x_15_n607), .ICO(M6_mult_x_15_n605), .CO(M6_mult_x_15_n606)
         );
  CMPR42X1 U26241 ( .A(M6_mult_x_15_n1100), .B(M6_mult_x_15_n1172), .C(
        M6_mult_x_15_n1148), .D(M6_mult_x_15_n648), .ICI(M6_mult_x_15_n1196), 
        .S(M6_mult_x_15_n640), .ICO(M6_mult_x_15_n638), .CO(M6_mult_x_15_n639)
         );
  CMPR42X1 U26242 ( .A(M6_mult_x_15_n652), .B(M6_mult_x_15_n1173), .C(
        M6_mult_x_15_n659), .D(M6_mult_x_15_n650), .ICI(M6_mult_x_15_n655), 
        .S(M6_mult_x_15_n647), .ICO(M6_mult_x_15_n645), .CO(M6_mult_x_15_n646)
         );
  CMPR42X1 U26243 ( .A(M6_mult_x_15_n1140), .B(M6_mult_x_15_n555), .C(
        M6_mult_x_15_n562), .D(M6_mult_x_15_n552), .ICI(M6_mult_x_15_n558), 
        .S(M6_mult_x_15_n549), .ICO(M6_mult_x_15_n547), .CO(M6_mult_x_15_n548)
         );
  CMPR42X1 U26244 ( .A(n22614), .B(n3220), .C(n10789), .D(M6_mult_x_15_n1017), 
        .ICI(M6_mult_x_15_n1064), .S(M6_mult_x_15_n515), .ICO(
        M6_mult_x_15_n513), .CO(M6_mult_x_15_n514) );
  CMPR42X1 U26245 ( .A(n26496), .B(n26494), .C(M6_mult_x_15_n1018), .D(
        M6_mult_x_15_n532), .ICI(M6_mult_x_15_n1041), .S(M6_mult_x_15_n524), 
        .ICO(M6_mult_x_15_n522), .CO(M6_mult_x_15_n523) );
  CMPR42X1 U26246 ( .A(M6_mult_x_15_n1165), .B(M6_mult_x_15_n1069), .C(
        M6_mult_x_15_n1117), .D(M6_mult_x_15_n1141), .ICI(M6_mult_x_15_n572), 
        .S(M6_mult_x_15_n563), .ICO(M6_mult_x_15_n561), .CO(M6_mult_x_15_n562)
         );
  CMPR42X1 U26247 ( .A(M6_mult_x_15_n567), .B(M6_mult_x_15_n557), .C(
        M6_mult_x_15_n1044), .D(M6_mult_x_15_n1164), .ICI(M6_mult_x_15_n561), 
        .S(M6_mult_x_15_n555), .ICO(M6_mult_x_15_n553), .CO(M6_mult_x_15_n554)
         );
  CMPR42X1 U26248 ( .A(M6_mult_x_15_n587), .B(M6_mult_x_15_n577), .C(
        M6_mult_x_15_n584), .D(M6_mult_x_15_n574), .ICI(M6_mult_x_15_n580), 
        .S(M6_mult_x_15_n571), .ICO(M6_mult_x_15_n569), .CO(M6_mult_x_15_n570)
         );
  CMPR42X1 U26249 ( .A(M6_mult_x_15_n1067), .B(M6_mult_x_15_n1139), .C(
        M6_mult_x_15_n553), .D(M6_mult_x_15_n550), .ICI(M6_mult_x_15_n554), 
        .S(M6_mult_x_15_n541), .ICO(M6_mult_x_15_n539), .CO(M6_mult_x_15_n540)
         );
  CMPR42X1 U26250 ( .A(M6_mult_x_15_n1102), .B(M6_mult_x_15_n1126), .C(
        M6_mult_x_15_n662), .D(M6_mult_x_15_n1174), .ICI(M6_mult_x_15_n668), 
        .S(M6_mult_x_15_n660), .ICO(M6_mult_x_15_n658), .CO(M6_mult_x_15_n659)
         );
  CMPR42X1 U26251 ( .A(M6_mult_x_15_n522), .B(M6_mult_x_15_n1040), .C(
        M6_mult_x_15_n1112), .D(M6_mult_x_15_n1088), .ICI(M6_mult_x_15_n523), 
        .S(M6_mult_x_15_n512), .ICO(M6_mult_x_15_n510), .CO(M6_mult_x_15_n511)
         );
  CMPR42X1 U26252 ( .A(M6_mult_x_15_n1061), .B(M6_mult_x_15_n492), .C(
        M6_mult_x_15_n486), .D(M6_mult_x_15_n493), .ICI(M6_mult_x_15_n489), 
        .S(M6_mult_x_15_n483), .ICO(M6_mult_x_15_n481), .CO(M6_mult_x_15_n482)
         );
  CMPR42X1 U26253 ( .A(M6_mult_x_15_n496), .B(M6_mult_x_15_n1062), .C(
        M6_mult_x_15_n502), .D(M6_mult_x_15_n494), .ICI(M6_mult_x_15_n498), 
        .S(M6_mult_x_15_n491), .ICO(M6_mult_x_15_n489), .CO(M6_mult_x_15_n490)
         );
  CMPR42X1 U26254 ( .A(M6_mult_x_15_n1060), .B(M6_mult_x_15_n484), .C(
        M6_mult_x_15_n479), .D(M6_mult_x_15_n485), .ICI(M6_mult_x_15_n481), 
        .S(M6_mult_x_15_n476), .ICO(M6_mult_x_15_n474), .CO(M6_mult_x_15_n475)
         );
  CMPR42X1 U26255 ( .A(M6_mult_x_15_n1035), .B(M6_mult_x_15_n1059), .C(
        M6_mult_x_15_n478), .D(M6_mult_x_15_n472), .ICI(M6_mult_x_15_n474), 
        .S(M6_mult_x_15_n469), .ICO(M6_mult_x_15_n467), .CO(M6_mult_x_15_n468)
         );
  CMPR42X1 U26256 ( .A(n22737), .B(n3217), .C(n11062), .D(M6_mult_x_15_n1011), 
        .ICI(M6_mult_x_15_n1058), .S(M6_mult_x_15_n466), .ICO(
        M6_mult_x_15_n464), .CO(M6_mult_x_15_n465) );
  CMPR42X1 U26257 ( .A(n26493), .B(n26491), .C(M6_mult_x_15_n1012), .D(
        M6_mult_x_15_n477), .ICI(M6_mult_x_15_n1083), .S(M6_mult_x_15_n472), 
        .ICO(M6_mult_x_15_n470), .CO(M6_mult_x_15_n471) );
  CMPR42X1 U26258 ( .A(n26489), .B(n9109), .C(n3219), .D(M6_mult_x_15_n1005), 
        .ICI(M6_mult_x_15_n436), .S(M6_mult_x_15_n435), .ICO(M6_mult_x_15_n433), .CO(M6_mult_x_15_n434) );
endmodule

